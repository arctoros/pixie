module Pixiez_Gamez_ofz_Life (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Not # (.UUID(64'd1173903214560679761 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_38), .out(wire_132));
  TC_Or3 # (.UUID(64'd3625327683154364378 ^ UUID), .BIT_WIDTH(64'd1)) Or3_1 (.in0(wire_320), .in1(wire_303), .in2(wire_250), .out(wire_88));
  TC_Or3 # (.UUID(64'd2550710310795524318 ^ UUID), .BIT_WIDTH(64'd1)) Or3_2 (.in0(wire_317), .in1(wire_269), .in2(wire_135), .out(wire_41));
  TC_Or3 # (.UUID(64'd2386266618142041082 ^ UUID), .BIT_WIDTH(64'd1)) Or3_3 (.in0(wire_380), .in1(wire_96), .in2(wire_81), .out(wire_436));
  TC_Or3 # (.UUID(64'd2492329720614052762 ^ UUID), .BIT_WIDTH(64'd1)) Or3_4 (.in0(wire_436), .in1(wire_41), .in2(wire_263), .out(wire_204));
  TC_Not # (.UUID(64'd798299516298535609 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_264), .out(wire_54));
  TC_DelayLine # (.UUID(64'd1033395116318490172 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_6 (.clk(clk), .rst(rst), .in(wire_54), .out(wire_264));
  TC_Not # (.UUID(64'd4512144033838034028 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_388), .out(wire_337));
  TC_Or3 # (.UUID(64'd3607001562755895464 ^ UUID), .BIT_WIDTH(64'd1)) Or3_8 (.in0(wire_108), .in1(wire_88), .in2(wire_130), .out(wire_388));
  TC_Add # (.UUID(64'd3899392937361653040 ^ UUID), .BIT_WIDTH(64'd8)) Add8_9 (.in0(wire_110), .in1(wire_251), .ci(wire_337), .out(wire_12), .co());
  TC_Or # (.UUID(64'd2898051740624681882 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_427), .in1(wire_266), .out(wire_320));
  TC_Not # (.UUID(64'd2990919190475442188 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_94), .out(wire_383));
  TC_Or3 # (.UUID(64'd275289339834281190 ^ UUID), .BIT_WIDTH(64'd1)) Or3_12 (.in0(wire_297), .in1(wire_175), .in2(wire_3), .out(wire_427));
  TC_Decoder3 # (.UUID(64'd4368521664392283939 ^ UUID)) Decoder3_13 (.dis(wire_360), .sel0(wire_57[0:0]), .sel1(wire_131[0:0]), .sel2(wire_56[0:0]), .out0(wire_317), .out1(wire_68), .out2(wire_29), .out3(wire_387), .out4(wire_11), .out5(wire_16), .out6(wire_3), .out7(wire_114));
  TC_Decoder3 # (.UUID(64'd2985802451890502143 ^ UUID)) Decoder3_14 (.dis(wire_174), .sel0(wire_57[0:0]), .sel1(wire_131[0:0]), .sel2(wire_56[0:0]), .out0(wire_220), .out1(wire_135), .out2(wire_269), .out3(wire_302), .out4(wire_193), .out5(wire_252), .out6(wire_156), .out7(wire_58));
  TC_Decoder3 # (.UUID(64'd3840069321658722899 ^ UUID)) Decoder3_15 (.dis(wire_283), .sel0(wire_57[0:0]), .sel1(wire_131[0:0]), .sel2(wire_56[0:0]), .out0(wire_243), .out1(wire_155), .out2(wire_42), .out3(wire_224), .out4(wire_61), .out5(wire_230), .out6(wire_127), .out7(wire_8));
  TC_Decoder3 # (.UUID(64'd2140688922873834327 ^ UUID)) Decoder3_16 (.dis(wire_373), .sel0(wire_57[0:0]), .sel1(wire_131[0:0]), .sel2(wire_56[0:0]), .out0(wire_183), .out1(wire_81), .out2(wire_96), .out3(wire_380), .out4(wire_100), .out5(wire_319), .out6(wire_119), .out7(wire_284));
  TC_Not # (.UUID(64'd2486164306052105983 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_434), .out(wire_360));
  TC_Not # (.UUID(64'd2538759475388196199 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_298), .out(wire_373));
  TC_Not # (.UUID(64'd2433569050415676182 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_205), .out(wire_283));
  TC_Not # (.UUID(64'd487282472206589942 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_342), .out(wire_174));
  TC_Maker8 # (.UUID(64'd3924075053356664533 ^ UUID)) Maker8_21 (.in0(wire_317), .in1(wire_68), .in2(wire_29), .in3(wire_387), .in4(wire_11), .in5(wire_16), .in6(wire_3), .in7(wire_114), .out(wire_165));
  TC_Maker8 # (.UUID(64'd4243729264906250734 ^ UUID)) Maker8_22 (.in0(wire_220), .in1(wire_135), .in2(wire_269), .in3(wire_302), .in4(wire_193), .in5(wire_252), .in6(wire_156), .in7(wire_58), .out(wire_141));
  TC_Maker8 # (.UUID(64'd3331907234886666019 ^ UUID)) Maker8_23 (.in0(wire_243), .in1(wire_155), .in2(wire_42), .in3(wire_224), .in4(wire_61), .in5(wire_230), .in6(wire_127), .in7(wire_8), .out(wire_189));
  TC_Maker8 # (.UUID(64'd1404105106470754509 ^ UUID)) Maker8_24 (.in0(wire_183), .in1(wire_81), .in2(wire_96), .in3(wire_380), .in4(wire_100), .in5(wire_319), .in6(wire_119), .in7(wire_284), .out(wire_288));
  TC_Or3 # (.UUID(64'd2149375025628133603 ^ UUID), .BIT_WIDTH(64'd1)) Or3_25 (.in0(wire_156), .in1(wire_58), .in2(wire_387), .out(wire_175));
  TC_Or3 # (.UUID(64'd3369381550219988481 ^ UUID), .BIT_WIDTH(64'd1)) Or3_26 (.in0(wire_319), .in1(wire_284), .in2(wire_243), .out(wire_266));
  TC_Or3 # (.UUID(64'd1730307490290969160 ^ UUID), .BIT_WIDTH(64'd1)) Or3_27 (.in0(wire_230), .in1(wire_61), .in2(wire_224), .out(wire_277));
  TC_Or3 # (.UUID(64'd1639935230616167963 ^ UUID), .BIT_WIDTH(64'd1)) Or3_28 (.in0(wire_220), .in1(wire_8), .in2(wire_127), .out(wire_365));
  TC_DelayLine # (.UUID(64'd4054610528999124272 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_29 (.clk(clk), .rst(rst), .in(wire_1[7:0]), .out(wire_109));
  TC_DelayLine # (.UUID(64'd4205670568223341846 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_209), .out(wire_38));
  TC_Splitter16 # (.UUID(64'd2407271182933992674 ^ UUID)) Splitter16_31 (.in(wire_187), .out0(wire_361), .out1(wire_191));
  TC_Maker16 # (.UUID(64'd3944115404361619184 ^ UUID)) Maker16_32 (.in0({{7{1'b0}}, wire_132 }), .in1(wire_394), .out(wire_187));
  TC_Or3 # (.UUID(64'd1442931798236221115 ^ UUID), .BIT_WIDTH(64'd1)) Or3_33 (.in0(wire_113), .in1(wire_43), .in2(wire_289), .out(wire_209));
  TC_Not # (.UUID(64'd610342714375567560 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_180[0:0]), .out(wire_435));
  TC_Not # (.UUID(64'd4450195243296613089 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_190[0:0]), .out(wire_201));
  TC_Splitter32 # (.UUID(64'd1978073918135016492 ^ UUID)) Splitter32_36 (.in(wire_170), .out0(wire_430), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd4139696140747098929 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_37 (.out(wire_423));
  TC_Mux # (.UUID(64'd4586296082639185111 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_14), .in0(wire_17), .in1(wire_423), .out(wire_356));
  TC_Add # (.UUID(64'd2939297397632065747 ^ UUID), .BIT_WIDTH(64'd8)) Add8_39 (.in0(wire_0), .in1(wire_356), .ci(1'd0), .out(wire_232), .co());
  TC_Mux # (.UUID(64'd4281127439128817208 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_40 (.sel(wire_133), .in0(wire_17), .in1(wire_307), .out(wire_393));
  TC_Neg # (.UUID(64'd2687713533780070524 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_41 (.in(wire_393), .out(wire_315));
  TC_Add # (.UUID(64'd594407689270678650 ^ UUID), .BIT_WIDTH(64'd8)) Add8_42 (.in0(wire_0), .in1(wire_315), .ci(1'd0), .out(wire_172), .co());
  TC_Mul # (.UUID(64'd3625573144411272462 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_43 (.in0(wire_0), .in1(wire_17), .out0(wire_177), .out1());
  TC_Switch # (.UUID(64'd924573676046716285 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_164), .in(wire_177), .out(wire_1_10[7:0]));
  TC_Switch # (.UUID(64'd3403135760287570862 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_267), .in(wire_172), .out(wire_1_15[7:0]));
  TC_Switch # (.UUID(64'd1563576092444781871 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_49), .in(wire_232), .out(wire_1_17[7:0]));
  TC_Splitter8 # (.UUID(64'd1279254792493053702 ^ UUID)) Splitter8_47 (.in(wire_430), .out0(wire_253), .out1(wire_310), .out2(wire_164), .out3(), .out4(wire_69), .out5(wire_14), .out6(wire_133), .out7(wire_35));
  TC_Not # (.UUID(64'd3866821846506759881 ^ UUID), .BIT_WIDTH(64'd1)) Not_48 (.in(wire_118[0:0]), .out(wire_329));
  TC_Switch # (.UUID(64'd2618318541541509822 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_94), .in(wire_160), .out(wire_0_1));
  TC_Switch # (.UUID(64'd4514760870899916219 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_383), .in(wire_160), .out(wire_255));
  TC_Switch # (.UUID(64'd92704038175830015 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_180[0:0]), .in(wire_186), .out(wire_17_0));
  TC_Switch # (.UUID(64'd3320542179656083506 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_435), .in(wire_186), .out(wire_182));
  TC_Switch # (.UUID(64'd2853649944201749510 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_118[0:0]), .in(wire_372), .out(wire_1_14[7:0]));
  TC_Switch # (.UUID(64'd1746760633635320209 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_329), .in(wire_372), .out(wire_281));
  TC_Splitter16 # (.UUID(64'd2696826286620571894 ^ UUID)) Splitter16_55 (.in(wire_323), .out0(wire_188), .out1(wire_190));
  TC_Or3 # (.UUID(64'd4510586934550576194 ^ UUID), .BIT_WIDTH(64'd1)) Or3_56 (.in0(wire_188[0:0]), .in1(wire_190[0:0]), .in2(wire_108), .out(wire_355));
  TC_Switch # (.UUID(64'd484565464453579756 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_188[0:0]), .in(wire_306[7:0]), .out(wire_291));
  TC_Switch # (.UUID(64'd2570328509294663425 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_58 (.en(wire_188[0:0]), .in(wire_45[7:0]), .out(wire_186));
  TC_Switch # (.UUID(64'd67298454145987374 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_59 (.en(wire_355), .in(wire_15[7:0]), .out(wire_160));
  TC_Mux # (.UUID(64'd2309406596842041848 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_60 (.sel(wire_201), .in0(wire_45[7:0]), .in1(wire_291), .out(wire_372));
  TC_Splitter16 # (.UUID(64'd3987227802858458071 ^ UUID)) Splitter16_61 (.in(wire_268), .out0(wire_118), .out1(wire_180));
  TC_Maker16 # (.UUID(64'd1122314457133455990 ^ UUID)) Maker16_62 (.in0({{7{1'b0}}, wire_413 }), .in1({{7{1'b0}}, wire_407 }), .out(wire_268));
  TC_Switch # (.UUID(64'd3625848211131814513 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_63 (.en(wire_38), .in(wire_109), .out(wire_394));
  TC_Mux # (.UUID(64'd2610902590828279325 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_64 (.sel(wire_361[0:0]), .in0(wire_191), .in1(wire_242), .out(wire_110));
  TC_Maker16 # (.UUID(64'd4154970328775153504 ^ UUID)) Maker16_65 (.in0({{7{1'b0}}, wire_130 }), .in1({{7{1'b0}}, wire_88 }), .out(wire_323));
  TC_Not # (.UUID(64'd1291016152359569471 ^ UUID), .BIT_WIDTH(64'd1)) Not_66 (.in(wire_54), .out(wire_218));
  TC_Counter # (.UUID(64'd4188127227668857882 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_67 (.clk(clk), .rst(rst), .save(wire_54), .in(wire_12), .out(wire_223));
  TC_Counter # (.UUID(64'd4007762735243366875 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_68 (.clk(clk), .rst(rst), .save(wire_264), .in(wire_12), .out(wire_438));
  TC_Switch # (.UUID(64'd1034539949200218368 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_69 (.en(wire_218), .in(wire_223), .out(wire_242_0));
  TC_Switch # (.UUID(64'd1470835681822839047 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_70 (.en(wire_54), .in(wire_438), .out(wire_242_1));
  TC_Constant # (.UUID(64'd4233708360558283991 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_71 (.out(wire_428));
  TC_Constant # (.UUID(64'd623194001325282984 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_72 (.out(wire_401));
  TC_Constant # (.UUID(64'd592794456182156764 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_73 (.out(wire_258));
  TC_Switch # (.UUID(64'd594207528242062231 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_74 (.en(wire_108), .in(wire_428), .out(wire_251_2));
  TC_Switch # (.UUID(64'd2669919813578549285 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_88), .in(wire_401), .out(wire_251_1));
  TC_Switch # (.UUID(64'd1342230075467448465 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_130), .in(wire_258), .out(wire_251_0));
  TC_Splitter8 # (.UUID(64'd335111286644642336 ^ UUID)) Splitter8_77 (.in(wire_31[7:0]), .out0(wire_71), .out1(wire_290), .out2(wire_326), .out3(wire_90), .out4(wire_139), .out5(wire_413), .out6(wire_407), .out7(wire_94));
  TC_Ram # (.UUID(64'd1796030558358045462 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_78 (.clk(clk), .rst(rst), .load(wire_40), .save(wire_22), .address({{24{1'b0}}, wire_198 }), .in0({{56{1'b0}}, wire_12 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_352), .out1(), .out2(), .out3());
  TC_Or # (.UUID(64'd1133444277294657592 ^ UUID), .BIT_WIDTH(64'd1)) Or_79 (.in0(wire_22), .in1(wire_40), .out(wire_113));
  TC_Splitter32 # (.UUID(64'd2085456252007348810 ^ UUID)) Splitter32_80 (.in(wire_170), .out0(), .out1(wire_10), .out2(), .out3(wire_158));
  TC_Or # (.UUID(64'd1885950073014372316 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_40), .in1(wire_22), .out(wire_378));
  TC_Switch # (.UUID(64'd3625428046281581986 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_82 (.en(wire_40), .in(wire_352[7:0]), .out(wire_1_19[7:0]));
  TC_Switch # (.UUID(64'd2958094378177111957 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_83 (.en(wire_22), .in(wire_0), .out(wire_1_18[7:0]));
  TC_Register # (.UUID(64'd188747501325143832 ^ UUID), .BIT_WIDTH(64'd8)) Register8_84 (.clk(clk), .rst(rst), .load(wire_378), .save(wire_378), .in(wire_363), .out(wire_93));
  TC_Switch # (.UUID(64'd412297402760837404 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_85 (.en(wire_22), .in(wire_424), .out(wire_363_0));
  TC_Switch # (.UUID(64'd2900436310909236685 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_86 (.en(wire_22), .in(wire_363), .out(wire_198_0));
  TC_Add # (.UUID(64'd257026951564140560 ^ UUID), .BIT_WIDTH(64'd8)) Add8_87 (.in0(wire_308), .in1(wire_93), .ci(1'd0), .out(wire_424), .co());
  TC_Switch # (.UUID(64'd1924045470845467746 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_88 (.en(wire_40), .in(wire_181), .out(wire_363_1));
  TC_Switch # (.UUID(64'd2699517944671878096 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_89 (.en(wire_40), .in(wire_93), .out(wire_198_1));
  TC_Constant # (.UUID(64'd114470560103204413 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_90 (.out(wire_308));
  TC_Neg # (.UUID(64'd1403767157571069852 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_91 (.in(wire_308), .out(wire_343));
  TC_Add # (.UUID(64'd226477113686883114 ^ UUID), .BIT_WIDTH(64'd8)) Add8_92 (.in0(wire_93), .in1(wire_343), .ci(1'd0), .out(wire_181), .co());
  TC_Constant # (.UUID(64'd1534915157065741767 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_93 (.out(wire_327));
  TC_Or # (.UUID(64'd250361279355801311 ^ UUID), .BIT_WIDTH(64'd1)) Or_94 (.in0(wire_92), .in1(wire_241), .out(wire_213));
  TC_LessU # (.UUID(64'd4052914289282609531 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_95 (.in0(wire_17), .in1(wire_0), .out(wire_241));
  TC_Not # (.UUID(64'd879017259160122171 ^ UUID), .BIT_WIDTH(64'd1)) Not_96 (.in(wire_92), .out(wire_325));
  TC_Or # (.UUID(64'd2827173067056184125 ^ UUID), .BIT_WIDTH(64'd1)) Or_97 (.in0(wire_227), .in1(wire_92), .out(wire_273));
  TC_Equal # (.UUID(64'd1702355244921692212 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_98 (.in0(wire_0), .in1(wire_17), .out(wire_92));
  TC_LessU # (.UUID(64'd2989501682613500020 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_99 (.in0(wire_0), .in1(wire_17), .out(wire_227));
  TC_Equal # (.UUID(64'd754200785245534088 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_100 (.in0(wire_327), .in1(wire_0), .out(wire_53));
  TC_Constant # (.UUID(64'd3349130739579016550 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_101 (.out(wire_154));
  TC_Switch # (.UUID(64'd4048450142757828966 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_102 (.en(wire_318), .in(wire_154), .out(wire_43_0));
  TC_Switch # (.UUID(64'd809238401857746034 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_103 (.en(wire_65), .in(wire_53), .out(wire_43_1));
  TC_Switch # (.UUID(64'd2006489762954213296 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_104 (.en(wire_64), .in(wire_227), .out(wire_43_2));
  TC_Switch # (.UUID(64'd3632517442940533649 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_105 (.en(wire_358), .in(wire_273), .out(wire_43_3));
  TC_Switch # (.UUID(64'd2587543755640527166 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_106 (.en(wire_221), .in(wire_92), .out(wire_43_4));
  TC_Switch # (.UUID(64'd4226160631432095931 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_107 (.en(wire_73), .in(wire_325), .out(wire_43_5));
  TC_Switch # (.UUID(64'd3303763842026803414 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_108 (.en(wire_261), .in(wire_213), .out(wire_43_6));
  TC_Switch # (.UUID(64'd2595133898896813930 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_109 (.en(wire_206), .in(wire_241), .out(wire_43_7));
  TC_Splitter8 # (.UUID(64'd4000441192049314171 ^ UUID)) Splitter8_110 (.in(wire_10), .out0(wire_318), .out1(wire_65), .out2(wire_64), .out3(wire_358), .out4(wire_221), .out5(wire_73), .out6(wire_261), .out7(wire_206));
  TC_Register # (.UUID(64'd1730520030450571584 ^ UUID), .BIT_WIDTH(64'd8)) Register8_111 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_399), .in(wire_1[7:0]), .out(wire_4));
  TC_Register # (.UUID(64'd2668217107469496786 ^ UUID), .BIT_WIDTH(64'd8)) Register8_112 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_212), .in(wire_1[7:0]), .out(wire_328));
  TC_Register # (.UUID(64'd3802042814775519440 ^ UUID), .BIT_WIDTH(64'd8)) Register8_113 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_126), .in(wire_1[7:0]), .out(wire_382));
  TC_Register # (.UUID(64'd3251616514511560897 ^ UUID), .BIT_WIDTH(64'd8)) Register8_114 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_9), .in(wire_1[7:0]), .out(wire_217));
  TC_Register # (.UUID(64'd3193651979249245240 ^ UUID), .BIT_WIDTH(64'd8)) Register8_115 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_162), .in(wire_1[7:0]), .out(wire_389));
  TC_Register # (.UUID(64'd3060613965044194374 ^ UUID), .BIT_WIDTH(64'd8)) Register8_116 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_333), .in(wire_1[7:0]), .out(wire_362));
  TC_Register # (.UUID(64'd323110644894396428 ^ UUID), .BIT_WIDTH(64'd8)) Register8_117 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_97), .in(wire_1[7:0]), .out(wire_28));
  TC_Register # (.UUID(64'd3914131157895841914 ^ UUID), .BIT_WIDTH(64'd8)) Register8_118 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_26), .in(wire_1[7:0]), .out(wire_366));
  TC_Register # (.UUID(64'd1377909213137338083 ^ UUID), .BIT_WIDTH(64'd8)) Register8_119 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_238), .in(wire_1[7:0]), .out(wire_331));
  TC_Register # (.UUID(64'd629828839776701115 ^ UUID), .BIT_WIDTH(64'd8)) Register8_120 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_321), .in(wire_1[7:0]), .out(wire_228));
  TC_Register # (.UUID(64'd3552817817526997674 ^ UUID), .BIT_WIDTH(64'd8)) Register8_121 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_305), .in(wire_1[7:0]), .out(wire_292));
  TC_Switch # (.UUID(64'd3583525001789596 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_122 (.en(wire_353), .in(wire_382), .out(wire_0_17));
  TC_Switch # (.UUID(64'd3589470201578893561 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_123 (.en(wire_19), .in(wire_382), .out(wire_17_16));
  TC_Switch # (.UUID(64'd3143479107291245555 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_124 (.en(wire_285), .in(wire_217), .out(wire_0_16));
  TC_Switch # (.UUID(64'd112316106613940142 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_125 (.en(wire_304), .in(wire_217), .out(wire_17_15));
  TC_Switch # (.UUID(64'd3379801696565704443 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_126 (.en(wire_121), .in(wire_28), .out(wire_0_15));
  TC_Switch # (.UUID(64'd2349617719032375395 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_127 (.en(wire_214), .in(wire_28), .out(wire_17_14));
  TC_Switch # (.UUID(64'd4345168894171961048 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_128 (.en(wire_87), .in(wire_331), .out(wire_0_14));
  TC_Switch # (.UUID(64'd1626712559099770596 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_129 (.en(wire_236), .in(wire_331), .out(wire_17_13));
  TC_Switch # (.UUID(64'd1791020341392350084 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_130 (.en(wire_322), .in(wire_366), .out(wire_0_13));
  TC_Switch # (.UUID(64'd2238730443596294210 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_131 (.en(wire_233), .in(wire_366), .out(wire_17_12));
  TC_Switch # (.UUID(64'd2319454654207709571 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_132 (.en(wire_364), .in(wire_389), .out(wire_0_12));
  TC_Switch # (.UUID(64'd3480139234004394235 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_133 (.en(wire_37), .in(wire_389), .out(wire_17_11));
  TC_Switch # (.UUID(64'd1188433479176944050 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_134 (.en(wire_46), .in(wire_228), .out(wire_0_11));
  TC_Switch # (.UUID(64'd1500034898745025292 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_135 (.en(wire_168), .in(wire_228), .out(wire_17_10));
  TC_Switch # (.UUID(64'd4328811457098718081 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_136 (.en(wire_210), .in(wire_362), .out(wire_0_10));
  TC_Switch # (.UUID(64'd2824054066706048507 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_137 (.en(wire_313), .in(wire_362), .out(wire_17_9));
  TC_Switch # (.UUID(64'd3566137095510004959 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_138 (.en(wire_13), .in(wire_328), .out(wire_0_9));
  TC_Switch # (.UUID(64'd1618994892661774692 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_139 (.en(wire_340), .in(wire_328), .out(wire_17_8));
  TC_Switch # (.UUID(64'd4518806407075154106 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_140 (.en(wire_301), .in(wire_4), .out(wire_0_8));
  TC_Switch # (.UUID(64'd4157847610664295546 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_141 (.en(wire_105), .in(wire_4), .out(wire_17_7));
  TC_Switch # (.UUID(64'd2520456579312250663 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_142 (.en(wire_62), .in(wire_292), .out(wire_0_7));
  TC_Switch # (.UUID(64'd891858636917436234 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_143 (.en(wire_178), .in(wire_292), .out(wire_17_6));
  TC_Switch # (.UUID(64'd1842801916941585222 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_144 (.en(wire_367), .in(wire_39), .out(wire_17_4));
  TC_Switch # (.UUID(64'd4332192567407784217 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_145 (.en(wire_256), .in(wire_39), .out(wire_0_5));
  TC_Switch # (.UUID(64'd2007288773695699471 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_146 (.en(wire_166), .in(wire_369), .out(wire_17_5));
  TC_Switch # (.UUID(64'd2659933361755871085 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_147 (.en(wire_246), .in(wire_369), .out(wire_0_6));
  TC_Register # (.UUID(64'd3909149542494051775 ^ UUID), .BIT_WIDTH(64'd8)) Register8_148 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_146), .in(wire_1[7:0]), .out(wire_369));
  TC_Register # (.UUID(64'd3813581101358275589 ^ UUID), .BIT_WIDTH(64'd8)) Register8_149 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_208), .in(wire_1[7:0]), .out(wire_39));
  TC_Splitter8 # (.UUID(64'd53967651305033637 ^ UUID)) Splitter8_150 (.in(wire_59), .out0(), .out1(), .out2(wire_34), .out3(wire_147), .out4(wire_22), .out5(wire_40), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd3641698352247847085 ^ UUID)) Splitter32_151 (.in(wire_170), .out0(), .out1(), .out2(), .out3(wire_59));
  TC_Switch # (.UUID(64'd3502727939898675348 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_152 (.en(wire_69), .in(wire_330), .out(wire_1_7[7:0]));
  TC_Switch # (.UUID(64'd3574082037932470167 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_153 (.en(wire_35), .in(wire_410), .out(wire_1_5[7:0]));
  TC_Neg # (.UUID(64'd2968407046620084969 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_154 (.in(wire_0), .out(wire_330));
  TC_Or # (.UUID(64'd2538623821936833797 ^ UUID), .BIT_WIDTH(64'd1)) Or_155 (.in0(wire_133), .in1(wire_310), .out(wire_267));
  TC_Constant # (.UUID(64'd1237391163366257378 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_156 (.out(wire_173));
  TC_Constant # (.UUID(64'd2599479896102896158 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_157 (.out(wire_307));
  TC_Ashr # (.UUID(64'd2161557586549500505 ^ UUID), .BIT_WIDTH(64'd8)) Ashr8_158 (.in(wire_0), .shift(wire_307), .out(wire_410));
  TC_Constant # (.UUID(64'd1556881997193880694 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_159 (.out(wire_24));
  TC_Switch # (.UUID(64'd3564139380929117312 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_160 (.en(wire_179), .in(wire_346), .out(wire_1_11[7:0]));
  TC_Switch # (.UUID(64'd111875663729447232 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_161 (.en(wire_104), .in(wire_23), .out(wire_1_8[7:0]));
  TC_And # (.UUID(64'd2752113776502556563 ^ UUID), .BIT_WIDTH(64'd8)) And8_162 (.in0(wire_0), .in1(wire_17), .out(wire_346));
  TC_Or # (.UUID(64'd1988259583830342258 ^ UUID), .BIT_WIDTH(64'd8)) Or8_163 (.in0(wire_0), .in1(wire_17), .out(wire_23));
  TC_Xor # (.UUID(64'd1084582658480022027 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_164 (.in0(wire_0), .in1(wire_17), .out(wire_21));
  TC_Not # (.UUID(64'd1474689859636581501 ^ UUID), .BIT_WIDTH(64'd8)) Not8_165 (.in(wire_0), .out(wire_390));
  TC_Shl # (.UUID(64'd1547575831449111006 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_166 (.in(wire_0), .shift(wire_173), .out(wire_144));
  TC_Shr # (.UUID(64'd120284355602086284 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_167 (.in(wire_0), .shift(wire_173), .out(wire_370));
  TC_Rol # (.UUID(64'd2716613345506561647 ^ UUID), .BIT_WIDTH(64'd8)) Rol8_168 (.in(wire_0), .shift(wire_173), .out(wire_137));
  TC_Ror # (.UUID(64'd1936902749111418424 ^ UUID), .BIT_WIDTH(64'd8)) Ror8_169 (.in(wire_0), .shift(wire_173), .out(wire_89));
  TC_Switch # (.UUID(64'd880910900980582870 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_170 (.en(wire_359), .in(wire_21), .out(wire_1_6[7:0]));
  TC_Switch # (.UUID(64'd3499157921667461283 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_171 (.en(wire_136), .in(wire_390), .out(wire_1_4[7:0]));
  TC_Switch # (.UUID(64'd2683242307298103541 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_172 (.en(wire_309), .in(wire_370), .out(wire_1_3[7:0]));
  TC_Switch # (.UUID(64'd2382702273644851040 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_173 (.en(wire_159), .in(wire_144), .out(wire_1_2[7:0]));
  TC_Switch # (.UUID(64'd3270310345322157611 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_174 (.en(wire_216), .in(wire_89), .out(wire_1_1[7:0]));
  TC_Switch # (.UUID(64'd2254212722512321080 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_175 (.en(wire_311), .in(wire_137), .out(wire_1_0[7:0]));
  TC_Splitter8 # (.UUID(64'd1804121337638409240 ^ UUID)) Splitter8_176 (.in(wire_6), .out0(wire_179), .out1(wire_104), .out2(wire_359), .out3(wire_136), .out4(wire_309), .out5(wire_159), .out6(wire_216), .out7(wire_311));
  TC_Splitter32 # (.UUID(64'd3827026339421898274 ^ UUID)) Splitter32_177 (.in(wire_170), .out0(), .out1(), .out2(wire_6), .out3());
  TC_Register # (.UUID(64'd2444082800644577615 ^ UUID), .BIT_WIDTH(64'd8)) Register8_178 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_237), .in(wire_1[7:0]), .out(wire_36));
  TC_Register # (.UUID(64'd2451162500981171780 ^ UUID), .BIT_WIDTH(64'd8)) Register8_179 (.clk(clk), .rst(rst), .load(wire_24), .save(wire_176), .in(wire_1[7:0]), .out(wire_271));
  TC_Switch # (.UUID(64'd4602360558464277168 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_180 (.en(wire_157), .in(wire_271), .out(wire_0_4));
  TC_Switch # (.UUID(64'd1030294617512356442 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_181 (.en(wire_50), .in(wire_271), .out(wire_17_3));
  TC_Switch # (.UUID(64'd3004960606798300169 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_182 (.en(wire_396), .in(wire_36), .out(wire_0_3));
  TC_Switch # (.UUID(64'd4002636313286681035 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_183 (.en(wire_229), .in(wire_36), .out(wire_17_2));
  TC_Switch # (.UUID(64'd1794948424895852344 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_184 (.en(wire_247), .in(wire_12), .out(wire_0_0));
  TC_Switch # (.UUID(64'd1973363098462495390 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_185 (.en(wire_125), .in(wire_12), .out(wire_17_1));
  TC_Or # (.UUID(64'd3685079247331042284 ^ UUID), .BIT_WIDTH(64'd1)) Or_186 (.in0(wire_98), .in1(wire_433), .out(wire_169));
  TC_Decoder3 # (.UUID(64'd1306852930812688709 ^ UUID)) Decoder3_187 (.dis(wire_254), .sel0(wire_91), .sel1(wire_134), .sel2(wire_260), .out0(wire_353), .out1(wire_285), .out2(wire_121), .out3(wire_87), .out4(wire_322), .out5(wire_364), .out6(wire_46), .out7(wire_210));
  TC_Decoder3 # (.UUID(64'd83913684500274929 ^ UUID)) Decoder3_188 (.dis(wire_169), .sel0(wire_91), .sel1(wire_134), .sel2(wire_260), .out0(wire_13), .out1(wire_301), .out2(wire_62), .out3(wire_246), .out4(wire_256), .out5(wire_157), .out6(wire_396), .out7());
  TC_Or # (.UUID(64'd77490688201718556 ^ UUID), .BIT_WIDTH(64'd1)) Or_189 (.in0(wire_106), .in1(wire_234), .out(wire_316));
  TC_Decoder3 # (.UUID(64'd1567803233114828732 ^ UUID)) Decoder3_190 (.dis(wire_257), .sel0(wire_75), .sel1(wire_129), .sel2(wire_138), .out0(wire_19), .out1(wire_304), .out2(wire_214), .out3(wire_236), .out4(wire_233), .out5(wire_37), .out6(wire_168), .out7(wire_313));
  TC_Decoder3 # (.UUID(64'd453336707101613734 ^ UUID)) Decoder3_191 (.dis(wire_316), .sel0(wire_75), .sel1(wire_129), .sel2(wire_138), .out0(wire_340), .out1(wire_105), .out2(wire_178), .out3(wire_166), .out4(wire_367), .out5(wire_50), .out6(wire_229), .out7());
  TC_Or # (.UUID(64'd3231982664529130647 ^ UUID), .BIT_WIDTH(64'd1)) Or_192 (.in0(wire_63), .in1(wire_194), .out(wire_376));
  TC_And # (.UUID(64'd1001988927217176368 ^ UUID), .BIT_WIDTH(64'd1)) And_193 (.in0(wire_30), .in1(wire_63), .out(wire_99));
  TC_Decoder3 # (.UUID(64'd881764854607920023 ^ UUID)) Decoder3_194 (.dis(wire_376), .sel0(wire_95), .sel1(wire_79), .sel2(wire_44), .out0(wire_212), .out1(wire_399), .out2(wire_305), .out3(wire_146), .out4(wire_208), .out5(wire_176), .out6(wire_237), .out7());
  TC_Decoder3 # (.UUID(64'd1290954479796467599 ^ UUID)) Decoder3_195 (.dis(wire_27), .sel0(wire_95), .sel1(wire_79), .sel2(wire_44), .out0(wire_126), .out1(wire_9), .out2(wire_97), .out3(wire_238), .out4(wire_26), .out5(wire_162), .out6(wire_321), .out7(wire_333));
  TC_Splitter8 # (.UUID(64'd836193493402382399 ^ UUID)) Splitter8_196 (.in(wire_281), .out0(wire_95), .out1(wire_79), .out2(wire_44), .out3(wire_30), .out4(wire_63), .out5(), .out6(), .out7());
  TC_Or3 # (.UUID(64'd1050286029460593336 ^ UUID), .BIT_WIDTH(64'd1)) Or3_197 (.in0(wire_365), .in1(wire_277), .in2(wire_425), .out(wire_263));
  TC_Or3 # (.UUID(64'd2135854994372188130 ^ UUID), .BIT_WIDTH(64'd1)) Or3_198 (.in0(wire_270[0:0]), .in1(wire_70), .in2(wire_106), .out(wire_257));
  TC_Not # (.UUID(64'd2526099756870330502 ^ UUID), .BIT_WIDTH(64'd1)) Not_199 (.in(wire_30), .out(wire_194));
  TC_Or3 # (.UUID(64'd2210994880038088801 ^ UUID), .BIT_WIDTH(64'd1)) Or3_200 (.in0(wire_351), .in1(wire_118[0:0]), .in2(wire_422), .out(wire_27));
  TC_Or3 # (.UUID(64'd2157493372619873439 ^ UUID), .BIT_WIDTH(64'd1)) Or3_201 (.in0(wire_249[0:0]), .in1(wire_52), .in2(wire_98), .out(wire_254));
  TC_And # (.UUID(64'd1226950749019374467 ^ UUID), .BIT_WIDTH(64'd1)) And_202 (.in0(wire_194), .in1(wire_63), .out(wire_289));
  TC_Splitter8 # (.UUID(64'd2422029773713477445 ^ UUID)) Splitter8_203 (.in(wire_182), .out0(wire_75), .out1(wire_129), .out2(wire_138), .out3(wire_70), .out4(wire_106), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd788460147325431136 ^ UUID), .BIT_WIDTH(64'd1)) And_204 (.in0(wire_106), .in1(wire_234), .out(wire_125));
  TC_Splitter8 # (.UUID(64'd3398032065560912619 ^ UUID)) Splitter8_205 (.in(wire_255), .out0(wire_91), .out1(wire_134), .out2(wire_260), .out3(wire_52), .out4(wire_98), .out5(), .out6(), .out7());
  TC_Maker32 # (.UUID(64'd4206831463159088388 ^ UUID)) Maker32_206 (.in0(wire_288), .in1(wire_189), .in2(wire_141), .in3(wire_165), .out(wire_170));
  TC_Or # (.UUID(64'd4008963988096052657 ^ UUID), .BIT_WIDTH(64'd1)) Or_207 (.in0(wire_14), .in1(wire_253), .out(wire_49));
  TC_Switch # (.UUID(64'd1437463996556091393 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_208 (.en(wire_278), .in(wire_0), .out(wire_1_12[7:0]));
  TC_Or3 # (.UUID(64'd4447495519109742911 ^ UUID), .BIT_WIDTH(64'd1)) Or3_209 (.in0(wire_29), .in1(wire_11), .in2(wire_16), .out(wire_108));
  TC_Or # (.UUID(64'd4073777860914098064 ^ UUID), .BIT_WIDTH(64'd1)) Or_210 (.in0(wire_11), .in1(wire_16), .out(wire_351));
  TC_Or # (.UUID(64'd3594630084656743215 ^ UUID), .BIT_WIDTH(64'd1)) Or_211 (.in0(wire_30), .in1(wire_63), .out(wire_422));
  TC_Splitter16 # (.UUID(64'd3981508339423121284 ^ UUID)) Splitter16_212 (.in(wire_196), .out0(wire_270), .out1(wire_249));
  TC_Maker16 # (.UUID(64'd905770393076995698 ^ UUID)) Maker16_213 (.in0(wire_180), .in1({{7{1'b0}}, wire_94 }), .out(wire_196));
  TC_Or3 # (.UUID(64'd3930544175131602979 ^ UUID), .BIT_WIDTH(64'd1)) Or3_214 (.in0(wire_302), .in1(wire_193), .in2(wire_252), .out(wire_297));
  TC_Program # (.UUID(64'd3486016637705709145 ^ UUID), .WORD_WIDTH(64'd32), .DEFAULT_FILE_NAME("Program_3060D1A98B8CE659.w32.bin"), .ARG_SIG("Program_3060D1A98B8CE659=%s")) Program_215 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_110 }), .out0(wire_31), .out1(wire_15), .out2(wire_45), .out3(wire_306));
  TC_Maker32 # (.UUID(64'd4293071912339536583 ^ UUID)) Maker32_216 (.in0({{7{1'b0}}, wire_71 }), .in1({{7{1'b0}}, wire_290 }), .in2({{7{1'b0}}, wire_326 }), .in3({{7{1'b0}}, wire_90 }), .out(wire_421));
  TC_Splitter32 # (.UUID(64'd1646892041393484876 ^ UUID)) Splitter32_217 (.in(wire_421), .out0(wire_57), .out1(wire_131), .out2(wire_56), .out3(wire_117));
  TC_Or # (.UUID(64'd431652671612996107 ^ UUID), .BIT_WIDTH(64'd1)) Or_218 (.in0(wire_119), .in1(wire_100), .out(wire_250));
  TC_Or # (.UUID(64'd3148152038805167791 ^ UUID), .BIT_WIDTH(64'd1)) Or_219 (.in0(wire_42), .in1(wire_183), .out(wire_425));
  TC_Or # (.UUID(64'd3136914901924744038 ^ UUID), .BIT_WIDTH(64'd1)) Or_220 (.in0(wire_68), .in1(wire_204), .out(wire_130));
  TC_Or # (.UUID(64'd915428529208528942 ^ UUID), .BIT_WIDTH(64'd1)) Or_221 (.in0(wire_155), .in1(wire_114), .out(wire_303));
  TC_Decoder2 # (.UUID(64'd586494721044460016 ^ UUID)) Decoder2_222 (.sel0(wire_117[0:0]), .sel1(wire_139), .out0(wire_298), .out1(wire_205), .out2(wire_342), .out3(wire_434));
  TC_Maker8 # (.UUID(64'd3779799189202718943 ^ UUID)) Maker8_223 (.in0(wire_349), .in1(wire_124), .in2(wire_374), .in3(wire_437), .in4(wire_344), .in5(wire_215), .in6(wire_350), .in7(wire_345), .out(wire_211));
  TC_Maker8 # (.UUID(64'd3170253293023823875 ^ UUID)) Maker8_224 (.in0(wire_240), .in1(wire_385), .in2(wire_414), .in3(wire_74), .in4(wire_225), .in5(wire_18), .in6(wire_426), .in7(wire_392), .out(wire_274));
  TC_Maker8 # (.UUID(64'd3132464070010384630 ^ UUID)) Maker8_225 (.in0(wire_391), .in1(wire_403), .in2(wire_280), .in3(wire_379), .in4(wire_419), .in5(wire_384), .in6(wire_219), .in7(wire_368), .out(wire_222));
  TC_Maker8 # (.UUID(64'd919537876160830977 ^ UUID)) Maker8_226 (.in0(wire_83), .in1(wire_336), .in2(wire_341), .in3(wire_192), .in4(wire_275), .in5(wire_185), .in6(wire_415), .in7(wire_357), .out(wire_420));
  TC_Maker8 # (.UUID(64'd977481532825068551 ^ UUID)) Maker8_227 (.in0(wire_397), .in1(wire_398), .in2(wire_416), .in3(wire_411), .in4(wire_202), .in5(wire_245), .in6(wire_279), .in7(wire_153), .out(wire_295));
  TC_Decoder3 # (.UUID(64'd2129725463425257505 ^ UUID)) Decoder3_228 (.dis(wire_171), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_349), .out1(wire_124), .out2(wire_374), .out3(wire_437), .out4(wire_344), .out5(wire_215), .out6(wire_350), .out7(wire_345));
  TC_Not # (.UUID(64'd3777762883375224886 ^ UUID), .BIT_WIDTH(64'd1)) Not_229 (.in(wire_76), .out(wire_123));
  TC_And # (.UUID(64'd4181286337335427174 ^ UUID), .BIT_WIDTH(64'd1)) And_230 (.in0(wire_347), .in1(wire_338), .out(wire_115));
  TC_And3 # (.UUID(64'd429931402316009848 ^ UUID), .BIT_WIDTH(64'd1)) And3_231 (.in0(wire_7), .in1(wire_248), .in2(wire_115), .out(wire_76));
  TC_And3 # (.UUID(64'd1928571948354264161 ^ UUID), .BIT_WIDTH(64'd1)) And3_232 (.in0(wire_207), .in1(wire_84), .in2(wire_78), .out(wire_140));
  TC_Not # (.UUID(64'd353608125405947400 ^ UUID), .BIT_WIDTH(64'd1)) Not_233 (.in(wire_84), .out(wire_248));
  TC_And3 # (.UUID(64'd3805392577439330749 ^ UUID), .BIT_WIDTH(64'd1)) And3_234 (.in0(wire_7), .in1(wire_148), .in2(wire_314), .out(wire_161));
  TC_And # (.UUID(64'd2972740437659232738 ^ UUID), .BIT_WIDTH(64'd1)) And_235 (.in0(wire_107), .in1(wire_395), .out(wire_314));
  TC_And3 # (.UUID(64'd1002689199071692242 ^ UUID), .BIT_WIDTH(64'd1)) And3_236 (.in0(wire_405), .in1(wire_417), .in2(wire_272), .out(wire_262));
  TC_And # (.UUID(64'd1231823558226297915 ^ UUID), .BIT_WIDTH(64'd1)) And_237 (.in0(wire_107), .in1(wire_282), .out(wire_272));
  TC_And3 # (.UUID(64'd2236749355694111481 ^ UUID), .BIT_WIDTH(64'd1)) And3_238 (.in0(wire_7), .in1(wire_84), .in2(wire_265), .out(wire_120));
  TC_And # (.UUID(64'd1468322473876195886 ^ UUID), .BIT_WIDTH(64'd1)) And_239 (.in0(wire_348), .in1(wire_101), .out(wire_265));
  TC_And # (.UUID(64'd4191888093249659745 ^ UUID), .BIT_WIDTH(64'd1)) And_240 (.in0(wire_259), .in1(wire_400), .out(wire_78));
  TC_Not # (.UUID(64'd4083524427655943283 ^ UUID), .BIT_WIDTH(64'd1)) Not_241 (.in(wire_85), .out(wire_395));
  TC_Not # (.UUID(64'd3079516046381206775 ^ UUID), .BIT_WIDTH(64'd1)) Not_242 (.in(wire_84), .out(wire_148));
  TC_Not # (.UUID(64'd3354472651210088626 ^ UUID), .BIT_WIDTH(64'd1)) Not_243 (.in(wire_7), .out(wire_405));
  TC_Not # (.UUID(64'd3736715756347921597 ^ UUID), .BIT_WIDTH(64'd1)) Not_244 (.in(wire_85), .out(wire_282));
  TC_Not # (.UUID(64'd114786921480515220 ^ UUID), .BIT_WIDTH(64'd1)) Not_245 (.in(wire_84), .out(wire_417));
  TC_Not # (.UUID(64'd226614187994715544 ^ UUID), .BIT_WIDTH(64'd1)) Not_246 (.in(wire_85), .out(wire_101));
  TC_Not # (.UUID(64'd99528564984418758 ^ UUID), .BIT_WIDTH(64'd1)) Not_247 (.in(wire_107), .out(wire_348));
  TC_Not # (.UUID(64'd3771918475425334235 ^ UUID), .BIT_WIDTH(64'd1)) Not_248 (.in(wire_7), .out(wire_207));
  TC_Not # (.UUID(64'd535351141032879899 ^ UUID), .BIT_WIDTH(64'd1)) Not_249 (.in(wire_85), .out(wire_400));
  TC_Not # (.UUID(64'd3324193097581102516 ^ UUID), .BIT_WIDTH(64'd1)) Not_250 (.in(wire_107), .out(wire_259));
  TC_Not # (.UUID(64'd195204682290887870 ^ UUID), .BIT_WIDTH(64'd1)) Not_251 (.in(wire_85), .out(wire_338));
  TC_Not # (.UUID(64'd1748957040376766845 ^ UUID), .BIT_WIDTH(64'd1)) Not_252 (.in(wire_107), .out(wire_347));
  TC_Not # (.UUID(64'd3967624677110085903 ^ UUID), .BIT_WIDTH(64'd1)) Not_253 (.in(wire_161), .out(wire_171));
  TC_Not # (.UUID(64'd275979249683281988 ^ UUID), .BIT_WIDTH(64'd1)) Not_254 (.in(wire_262), .out(wire_432));
  TC_Not # (.UUID(64'd3166221433695873745 ^ UUID), .BIT_WIDTH(64'd1)) Not_255 (.in(wire_120), .out(wire_197));
  TC_Not # (.UUID(64'd2659467157919984791 ^ UUID), .BIT_WIDTH(64'd1)) Not_256 (.in(wire_140), .out(wire_111));
  TC_Splitter8 # (.UUID(64'd305375785571403410 ^ UUID)) Splitter8_257 (.in(wire_112), .out0(wire_60), .out1(wire_25), .out2(wire_5), .out3(wire_7), .out4(wire_84), .out5(wire_107), .out6(wire_85), .out7());
  TC_Decoder3 # (.UUID(64'd2111100196510366165 ^ UUID)) Decoder3_258 (.dis(wire_432), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_240), .out1(wire_385), .out2(wire_414), .out3(wire_74), .out4(wire_225), .out5(wire_18), .out6(wire_426), .out7(wire_392));
  TC_Decoder3 # (.UUID(64'd3300166719084188568 ^ UUID)) Decoder3_259 (.dis(wire_197), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_391), .out1(wire_403), .out2(wire_280), .out3(wire_379), .out4(wire_419), .out5(wire_384), .out6(wire_219), .out7(wire_368));
  TC_Decoder3 # (.UUID(64'd3552639083627078804 ^ UUID)) Decoder3_260 (.dis(wire_111), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_83), .out1(wire_336), .out2(wire_341), .out3(wire_192), .out4(wire_275), .out5(wire_185), .out6(wire_415), .out7(wire_357));
  TC_Decoder3 # (.UUID(64'd720807239010054970 ^ UUID)) Decoder3_261 (.dis(wire_123), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_397), .out1(wire_398), .out2(wire_416), .out3(wire_411), .out4(wire_202), .out5(wire_245), .out6(wire_279), .out7(wire_153));
  TC_Maker8 # (.UUID(64'd580009802560296023 ^ UUID)) Maker8_262 (.in0(wire_48), .in1(wire_163), .in2(wire_276), .in3(wire_32), .in4(wire_339), .in5(wire_299), .in6(wire_402), .in7(wire_312), .out(wire_116));
  TC_Not # (.UUID(64'd1034141622614219055 ^ UUID), .BIT_WIDTH(64'd1)) Not_263 (.in(wire_107), .out(wire_404));
  TC_Not # (.UUID(64'd4484983783826623864 ^ UUID), .BIT_WIDTH(64'd1)) Not_264 (.in(wire_85), .out(wire_184));
  TC_Decoder3 # (.UUID(64'd4451693059702490902 ^ UUID)) Decoder3_265 (.dis(wire_231), .sel0(wire_60), .sel1(wire_25), .sel2(wire_5), .out0(wire_48), .out1(wire_163), .out2(wire_276), .out3(wire_32), .out4(wire_339), .out5(wire_299), .out6(wire_402), .out7(wire_312));
  TC_And3 # (.UUID(64'd345998752798203089 ^ UUID), .BIT_WIDTH(64'd1)) And3_266 (.in0(wire_99), .in1(wire_404), .in2(wire_184), .out(wire_226));
  TC_Add # (.UUID(64'd2292127294728674804 ^ UUID), .BIT_WIDTH(64'd8)) Add8_267 (.in0(wire_122), .in1(wire_20), .ci(1'd0), .out(wire_112), .co());
  TC_Constant # (.UUID(64'd3974248596445317617 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_268 (.out(wire_72));
  TC_Not # (.UUID(64'd3228970102034108709 ^ UUID), .BIT_WIDTH(64'd1)) Not_269 (.in(wire_7), .out(wire_287));
  TC_Not # (.UUID(64'd4020811955063250824 ^ UUID), .BIT_WIDTH(64'd1)) Not_270 (.in(wire_84), .out(wire_77));
  TC_Not # (.UUID(64'd3082843848025648527 ^ UUID), .BIT_WIDTH(64'd1)) Not_271 (.in(wire_145), .out(wire_231));
  TC_And3 # (.UUID(64'd1984641945363423930 ^ UUID), .BIT_WIDTH(64'd1)) And3_272 (.in0(wire_287), .in1(wire_77), .in2(wire_226), .out(wire_145));
  TC_And # (.UUID(64'd1124549664905356862 ^ UUID), .BIT_WIDTH(64'd8)) And8_273 (.in0(wire_150), .in1(wire_151), .out(wire_20));
  TC_Constant # (.UUID(64'd985218960685118192 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h60)) Constant8_274 (.out(wire_408));
  TC_Constant # (.UUID(64'd261774725404830716 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h30)) Constant8_275 (.out(wire_128));
  TC_Neg # (.UUID(64'd4080209337533804453 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_276 (.in(wire_167), .out(wire_122));
  TC_Switch # (.UUID(64'd1589832099590329381 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_277 (.en(wire_244), .in(wire_408), .out(wire_167_0));
  TC_Switch # (.UUID(64'd3370031454424542084 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_278 (.en(wire_67), .in(wire_128), .out(wire_167_1));
  TC_DotMatrixDisplay # (.UUID(64'd4414540759399644336 ^ UUID)) DotMatrixDisplay_279 (.clk(clk), .rst(rst), .en_y(wire_293[0:0]), .en_x(wire_102[0:0]), .color_info(wire_293), .pixel_info(wire_102));
  TC_DotMatrixDisplay # (.UUID(64'd1220696841797878838 ^ UUID)) DotMatrixDisplay_280 (.clk(clk), .rst(rst), .en_y(wire_200[0:0]), .en_x(wire_102[0:0]), .color_info(wire_200), .pixel_info(wire_102));
  TC_DotMatrixDisplay # (.UUID(64'd2805810588850820154 ^ UUID)) DotMatrixDisplay_281 (.clk(clk), .rst(rst), .en_y(wire_286[0:0]), .en_x(wire_102[0:0]), .color_info(wire_286), .pixel_info(wire_102));
  TC_Constant # (.UUID(64'd3274466395144906983 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h30)) Constant8_282 (.out(wire_418));
  TC_Maker32 # (.UUID(64'd1996266684949409194 ^ UUID)) Maker32_283 (.in0({{7{1'b0}}, wire_67 }), .in1(wire_429), .in2(wire_354), .in3(wire_371), .out(wire_200));
  TC_LessU # (.UUID(64'd2002074936609615378 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_284 (.in0(wire_20), .in1(wire_334), .out(wire_103));
  TC_LessU # (.UUID(64'd862924152651395411 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_285 (.in0(wire_20), .in1(wire_386), .out(wire_377));
  TC_LessU # (.UUID(64'd2376808415796356142 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_286 (.in0(wire_20), .in1(wire_418), .out(wire_51));
  TC_Constant # (.UUID(64'd1564012343140950201 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h80)) Constant8_287 (.out(wire_334));
  TC_Constant # (.UUID(64'd3863067129706704118 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h60)) Constant8_288 (.out(wire_386));
  TC_Not # (.UUID(64'd573075325026521668 ^ UUID), .BIT_WIDTH(64'd1)) Not_289 (.in(wire_377), .out(wire_82));
  TC_Not # (.UUID(64'd481913933217625022 ^ UUID), .BIT_WIDTH(64'd1)) Not_290 (.in(wire_51), .out(wire_381));
  TC_Not # (.UUID(64'd4550021201972865238 ^ UUID), .BIT_WIDTH(64'd1)) Not_291 (.in(wire_51), .out(wire_86));
  TC_And3 # (.UUID(64'd748936417975850292 ^ UUID), .BIT_WIDTH(64'd1)) And3_292 (.in0(wire_381), .in1(wire_82), .in2(wire_103), .out(wire_244));
  TC_And3 # (.UUID(64'd2074191732282209651 ^ UUID), .BIT_WIDTH(64'd1)) And3_293 (.in0(wire_86), .in1(wire_377), .in2(wire_103), .out(wire_67));
  TC_And3 # (.UUID(64'd1126180895750929946 ^ UUID), .BIT_WIDTH(64'd1)) And3_294 (.in0(wire_51), .in1(wire_377), .in2(wire_103), .out(wire_239));
  TC_Maker64 # (.UUID(64'd1315198523453947527 ^ UUID)) Maker64_295 (.in0({{7{1'b0}}, wire_72 }), .in1(wire_116), .in2(wire_295), .in3(wire_420), .in4(wire_222), .in5(wire_274), .in6(wire_211), .in7({{7{1'b0}}, wire_72 }), .out(wire_102));
  TC_Maker32 # (.UUID(64'd4008862029770199109 ^ UUID)) Maker32_296 (.in0({{7{1'b0}}, wire_244 }), .in1(wire_235), .in2(wire_142), .in3(wire_375), .out(wire_286));
  TC_Maker32 # (.UUID(64'd1250450978058653133 ^ UUID)) Maker32_297 (.in0({{7{1'b0}}, wire_239 }), .in1(wire_195), .in2(wire_324), .in3(wire_406), .out(wire_293));
  TC_Splitter32 # (.UUID(64'd4207847732869802758 ^ UUID)) Splitter32_298 (.in(wire_66), .out0(), .out1(wire_195), .out2(wire_324), .out3(wire_406));
  TC_Splitter32 # (.UUID(64'd1250593027688444578 ^ UUID)) Splitter32_299 (.in(wire_66), .out0(), .out1(wire_429), .out2(wire_354), .out3(wire_371));
  TC_Splitter32 # (.UUID(64'd174210753003038335 ^ UUID)) Splitter32_300 (.in(wire_66), .out0(), .out1(wire_235), .out2(wire_142), .out3(wire_375));
  TC_LessU # (.UUID(64'd362456343450182185 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_301 (.in0(wire_150), .in1(wire_151), .out(wire_332));
  TC_Constant # (.UUID(64'd712959216000692405 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7F)) Constant8_302 (.out(wire_150));
  TC_Constant # (.UUID(64'd2673145422975682581 ^ UUID), .BIT_WIDTH(64'd32), .value(32'hFFFFFF00)) Constant32_303 (.out(wire_296));
  TC_Switch # (.UUID(64'd521043265076875738 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_304 (.en(wire_332), .in(wire_296), .out(wire_66));
  TC_Not # (.UUID(64'd650880247707744954 ^ UUID), .BIT_WIDTH(64'd1)) Not_305 (.in(wire_70), .out(wire_234));
  TC_Ram # (.UUID(64'd4026031931514975637 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_306 (.clk(clk), .rst(rst), .load(wire_147), .save(wire_34), .address({{24{1'b0}}, wire_55 }), .in0({{56{1'b0}}, wire_0 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_1_9), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd3186469103346041057 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_307 (.out(wire_335));
  TC_Neg # (.UUID(64'd1596347693989418526 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_308 (.in(wire_335), .out(wire_409));
  TC_Register # (.UUID(64'd3208768588500146265 ^ UUID), .BIT_WIDTH(64'd8)) Register8_309 (.clk(clk), .rst(rst), .load(wire_203), .save(wire_203), .in(wire_199), .out(wire_47));
  TC_Switch # (.UUID(64'd2570549170391169806 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_310 (.en(wire_34), .in(wire_412), .out(wire_199_0));
  TC_Switch # (.UUID(64'd1292048990515190170 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_311 (.en(wire_34), .in(wire_199), .out(wire_55_0));
  TC_Add # (.UUID(64'd64358517018617917 ^ UUID), .BIT_WIDTH(64'd8)) Add8_312 (.in0(wire_335), .in1(wire_47), .ci(1'd0), .out(wire_412), .co());
  TC_Switch # (.UUID(64'd1472851788000812976 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_313 (.en(wire_147), .in(wire_149), .out(wire_199_1));
  TC_Switch # (.UUID(64'd3926632308267132297 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_314 (.en(wire_147), .in(wire_47), .out(wire_55_1));
  TC_Or # (.UUID(64'd3243870362582900008 ^ UUID), .BIT_WIDTH(64'd1)) Or_315 (.in0(wire_147), .in1(wire_34), .out(wire_203));
  TC_Add # (.UUID(64'd901104549422042229 ^ UUID), .BIT_WIDTH(64'd8)) Add8_316 (.in0(wire_47), .in1(wire_409), .ci(1'd0), .out(wire_149), .co());
  TC_Ram # (.UUID(64'd1246387032842321975 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_317 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_143), .address({{24{1'b0}}, wire_17 }), .in0({{56{1'b0}}, wire_0 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_1_16), .out1(), .out2(), .out3());
  TC_Splitter8 # (.UUID(64'd4075614425899748182 ^ UUID)) Splitter8_318 (.in(wire_158), .out0(wire_143), .out1(wire_2), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_278));
  TC_Program # (.UUID(64'd2888906506993602274 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_281775297AAB0EE2.w8.bin"), .ARG_SIG("Program_281775297AAB0EE2=%s")) Program_319 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_0 }), .out0(wire_152), .out1(), .out2(), .out3());
  TC_Switch # (.UUID(64'd2910385312128859062 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_320 (.en(wire_33), .in(wire_152[7:0]), .out(wire_1_13[7:0]));
  TC_Timing # (.UUID(64'd213808295465521726 ^ UUID)) Timing_321 (.en(wire_431), .out(wire_300));
  TC_Constant # (.UUID(64'd4167380902895038125 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_322 (.out(wire_431));
  TC_Splitter8 # (.UUID(64'd321008928267196602 ^ UUID)) Splitter8_323 (.in(wire_288), .out0(), .out1(), .out2(), .out3(wire_33), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd2205580488541737701 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_324 (.en(wire_80), .in(wire_300[0:0]), .out(wire_0_2[0:0]));
  TC_Not # (.UUID(64'd4572459903145988353 ^ UUID), .BIT_WIDTH(64'd1)) Not_325 (.in(wire_52), .out(wire_433));
  TC_And # (.UUID(64'd2959708723279158992 ^ UUID), .BIT_WIDTH(64'd1)) And_326 (.in0(wire_52), .in1(wire_98), .out(wire_80));
  TC_And # (.UUID(64'd2938706705872922893 ^ UUID), .BIT_WIDTH(64'd1)) And_327 (.in0(wire_98), .in1(wire_294), .out(wire_247));
  TC_Not # (.UUID(64'd2047231847930482224 ^ UUID), .BIT_WIDTH(64'd1)) Not_328 (.in(wire_52), .out(wire_294));
  TC_Switch # (.UUID(64'd1215961827164946147 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_329 (.en(wire_99), .in(wire_1[7:0]), .out(wire_151));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  wire [7:0] wire_0_4;
  wire [7:0] wire_0_5;
  wire [7:0] wire_0_6;
  wire [7:0] wire_0_7;
  wire [7:0] wire_0_8;
  wire [7:0] wire_0_9;
  wire [7:0] wire_0_10;
  wire [7:0] wire_0_11;
  wire [7:0] wire_0_12;
  wire [7:0] wire_0_13;
  wire [7:0] wire_0_14;
  wire [7:0] wire_0_15;
  wire [7:0] wire_0_16;
  wire [7:0] wire_0_17;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6|wire_0_7|wire_0_8|wire_0_9|wire_0_10|wire_0_11|wire_0_12|wire_0_13|wire_0_14|wire_0_15|wire_0_16|wire_0_17;
  wire [63:0] wire_1;
  wire [63:0] wire_1_0;
  wire [63:0] wire_1_1;
  wire [63:0] wire_1_2;
  wire [63:0] wire_1_3;
  wire [63:0] wire_1_4;
  wire [63:0] wire_1_5;
  wire [63:0] wire_1_6;
  wire [63:0] wire_1_7;
  wire [63:0] wire_1_8;
  wire [63:0] wire_1_9;
  wire [63:0] wire_1_10;
  wire [63:0] wire_1_11;
  wire [63:0] wire_1_12;
  wire [63:0] wire_1_13;
  wire [63:0] wire_1_14;
  wire [63:0] wire_1_15;
  wire [63:0] wire_1_16;
  wire [63:0] wire_1_17;
  wire [63:0] wire_1_18;
  wire [63:0] wire_1_19;
  assign wire_1 = wire_1_0|wire_1_1|wire_1_2|wire_1_3|wire_1_4|wire_1_5|wire_1_6|wire_1_7|wire_1_8|wire_1_9|wire_1_10|wire_1_11|wire_1_12|wire_1_13|wire_1_14|wire_1_15|wire_1_16|wire_1_17|wire_1_18|wire_1_19;
  wire [0:0] wire_2;
  wire [0:0] wire_3;
  wire [7:0] wire_4;
  wire [0:0] wire_5;
  wire [7:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [0:0] wire_13;
  wire [0:0] wire_14;
  wire [63:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [7:0] wire_17_0;
  wire [7:0] wire_17_1;
  wire [7:0] wire_17_2;
  wire [7:0] wire_17_3;
  wire [7:0] wire_17_4;
  wire [7:0] wire_17_5;
  wire [7:0] wire_17_6;
  wire [7:0] wire_17_7;
  wire [7:0] wire_17_8;
  wire [7:0] wire_17_9;
  wire [7:0] wire_17_10;
  wire [7:0] wire_17_11;
  wire [7:0] wire_17_12;
  wire [7:0] wire_17_13;
  wire [7:0] wire_17_14;
  wire [7:0] wire_17_15;
  wire [7:0] wire_17_16;
  assign wire_17 = wire_17_0|wire_17_1|wire_17_2|wire_17_3|wire_17_4|wire_17_5|wire_17_6|wire_17_7|wire_17_8|wire_17_9|wire_17_10|wire_17_11|wire_17_12|wire_17_13|wire_17_14|wire_17_15|wire_17_16;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [7:0] wire_21;
  wire [0:0] wire_22;
  wire [7:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [7:0] wire_28;
  wire [0:0] wire_29;
  wire [0:0] wire_30;
  wire [63:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [7:0] wire_36;
  wire [0:0] wire_37;
  wire [0:0] wire_38;
  wire [7:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [0:0] wire_43_0;
  wire [0:0] wire_43_1;
  wire [0:0] wire_43_2;
  wire [0:0] wire_43_3;
  wire [0:0] wire_43_4;
  wire [0:0] wire_43_5;
  wire [0:0] wire_43_6;
  wire [0:0] wire_43_7;
  assign wire_43 = wire_43_0|wire_43_1|wire_43_2|wire_43_3|wire_43_4|wire_43_5|wire_43_6|wire_43_7;
  wire [0:0] wire_44;
  wire [63:0] wire_45;
  wire [0:0] wire_46;
  wire [7:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [7:0] wire_55_0;
  wire [7:0] wire_55_1;
  assign wire_55 = wire_55_0|wire_55_1;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [7:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [0:0] wire_62;
  wire [0:0] wire_63;
  wire [0:0] wire_64;
  wire [0:0] wire_65;
  wire [31:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [0:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [0:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [7:0] wire_89;
  wire [0:0] wire_90;
  wire [0:0] wire_91;
  wire [0:0] wire_92;
  wire [7:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [63:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [7:0] wire_109;
  wire [7:0] wire_110;
  wire [0:0] wire_111;
  wire [7:0] wire_112;
  wire [0:0] wire_113;
  wire [0:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [7:0] wire_117;
  wire [7:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [7:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;
  wire [0:0] wire_127;
  wire [7:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [7:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [0:0] wire_135;
  wire [0:0] wire_136;
  wire [7:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [7:0] wire_141;
  wire [7:0] wire_142;
  wire [0:0] wire_143;
  wire [7:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [0:0] wire_147;
  wire [0:0] wire_148;
  wire [7:0] wire_149;
  wire [7:0] wire_150;
  wire [7:0] wire_151;
  wire [63:0] wire_152;
  wire [0:0] wire_153;
  wire [0:0] wire_154;
  wire [0:0] wire_155;
  wire [0:0] wire_156;
  wire [0:0] wire_157;
  wire [7:0] wire_158;
  wire [0:0] wire_159;
  wire [7:0] wire_160;
  wire [0:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [7:0] wire_165;
  wire [0:0] wire_166;
  wire [7:0] wire_167;
  wire [7:0] wire_167_0;
  wire [7:0] wire_167_1;
  assign wire_167 = wire_167_0|wire_167_1;
  wire [0:0] wire_168;
  wire [0:0] wire_169;
  wire [31:0] wire_170;
  wire [0:0] wire_171;
  wire [7:0] wire_172;
  wire [7:0] wire_173;
  wire [0:0] wire_174;
  wire [0:0] wire_175;
  wire [0:0] wire_176;
  wire [7:0] wire_177;
  wire [0:0] wire_178;
  wire [0:0] wire_179;
  wire [7:0] wire_180;
  wire [7:0] wire_181;
  wire [7:0] wire_182;
  wire [0:0] wire_183;
  wire [0:0] wire_184;
  wire [0:0] wire_185;
  wire [7:0] wire_186;
  wire [15:0] wire_187;
  wire [7:0] wire_188;
  wire [7:0] wire_189;
  wire [7:0] wire_190;
  wire [7:0] wire_191;
  wire [0:0] wire_192;
  wire [0:0] wire_193;
  wire [0:0] wire_194;
  wire [7:0] wire_195;
  wire [15:0] wire_196;
  wire [0:0] wire_197;
  wire [7:0] wire_198;
  wire [7:0] wire_198_0;
  wire [7:0] wire_198_1;
  assign wire_198 = wire_198_0|wire_198_1;
  wire [7:0] wire_199;
  wire [7:0] wire_199_0;
  wire [7:0] wire_199_1;
  assign wire_199 = wire_199_0|wire_199_1;
  wire [31:0] wire_200;
  wire [0:0] wire_201;
  wire [0:0] wire_202;
  wire [0:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [0:0] wire_206;
  wire [0:0] wire_207;
  wire [0:0] wire_208;
  wire [0:0] wire_209;
  wire [0:0] wire_210;
  wire [7:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [0:0] wire_214;
  wire [0:0] wire_215;
  wire [0:0] wire_216;
  wire [7:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [0:0] wire_221;
  wire [7:0] wire_222;
  wire [7:0] wire_223;
  wire [0:0] wire_224;
  wire [0:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [7:0] wire_228;
  wire [0:0] wire_229;
  wire [0:0] wire_230;
  wire [0:0] wire_231;
  wire [7:0] wire_232;
  wire [0:0] wire_233;
  wire [0:0] wire_234;
  wire [7:0] wire_235;
  wire [0:0] wire_236;
  wire [0:0] wire_237;
  wire [0:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [7:0] wire_242;
  wire [7:0] wire_242_0;
  wire [7:0] wire_242_1;
  assign wire_242 = wire_242_0|wire_242_1;
  wire [0:0] wire_243;
  wire [0:0] wire_244;
  wire [0:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [0:0] wire_248;
  wire [7:0] wire_249;
  wire [0:0] wire_250;
  wire [7:0] wire_251;
  wire [7:0] wire_251_0;
  wire [7:0] wire_251_1;
  wire [7:0] wire_251_2;
  assign wire_251 = wire_251_0|wire_251_1|wire_251_2;
  wire [0:0] wire_252;
  wire [0:0] wire_253;
  wire [0:0] wire_254;
  wire [7:0] wire_255;
  wire [0:0] wire_256;
  wire [0:0] wire_257;
  wire [7:0] wire_258;
  wire [0:0] wire_259;
  wire [0:0] wire_260;
  wire [0:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [0:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [15:0] wire_268;
  wire [0:0] wire_269;
  wire [7:0] wire_270;
  wire [7:0] wire_271;
  wire [0:0] wire_272;
  wire [0:0] wire_273;
  wire [7:0] wire_274;
  wire [0:0] wire_275;
  wire [0:0] wire_276;
  wire [0:0] wire_277;
  wire [0:0] wire_278;
  wire [0:0] wire_279;
  wire [0:0] wire_280;
  wire [7:0] wire_281;
  wire [0:0] wire_282;
  wire [0:0] wire_283;
  wire [0:0] wire_284;
  wire [0:0] wire_285;
  wire [31:0] wire_286;
  wire [0:0] wire_287;
  wire [7:0] wire_288;
  wire [0:0] wire_289;
  wire [0:0] wire_290;
  wire [7:0] wire_291;
  wire [7:0] wire_292;
  wire [31:0] wire_293;
  wire [0:0] wire_294;
  wire [7:0] wire_295;
  wire [31:0] wire_296;
  wire [0:0] wire_297;
  wire [0:0] wire_298;
  wire [0:0] wire_299;
  wire [63:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [0:0] wire_303;
  wire [0:0] wire_304;
  wire [0:0] wire_305;
  wire [63:0] wire_306;
  wire [7:0] wire_307;
  wire [7:0] wire_308;
  wire [0:0] wire_309;
  wire [0:0] wire_310;
  wire [0:0] wire_311;
  wire [0:0] wire_312;
  wire [0:0] wire_313;
  wire [0:0] wire_314;
  wire [7:0] wire_315;
  wire [0:0] wire_316;
  wire [0:0] wire_317;
  wire [0:0] wire_318;
  wire [0:0] wire_319;
  wire [0:0] wire_320;
  wire [0:0] wire_321;
  wire [0:0] wire_322;
  wire [15:0] wire_323;
  wire [7:0] wire_324;
  wire [0:0] wire_325;
  wire [0:0] wire_326;
  wire [7:0] wire_327;
  wire [7:0] wire_328;
  wire [0:0] wire_329;
  wire [7:0] wire_330;
  wire [7:0] wire_331;
  wire [0:0] wire_332;
  wire [0:0] wire_333;
  wire [7:0] wire_334;
  wire [7:0] wire_335;
  wire [0:0] wire_336;
  wire [0:0] wire_337;
  wire [0:0] wire_338;
  wire [0:0] wire_339;
  wire [0:0] wire_340;
  wire [0:0] wire_341;
  wire [0:0] wire_342;
  wire [7:0] wire_343;
  wire [0:0] wire_344;
  wire [0:0] wire_345;
  wire [7:0] wire_346;
  wire [0:0] wire_347;
  wire [0:0] wire_348;
  wire [0:0] wire_349;
  wire [0:0] wire_350;
  wire [0:0] wire_351;
  wire [63:0] wire_352;
  wire [0:0] wire_353;
  wire [7:0] wire_354;
  wire [0:0] wire_355;
  wire [7:0] wire_356;
  wire [0:0] wire_357;
  wire [0:0] wire_358;
  wire [0:0] wire_359;
  wire [0:0] wire_360;
  wire [7:0] wire_361;
  wire [7:0] wire_362;
  wire [7:0] wire_363;
  wire [7:0] wire_363_0;
  wire [7:0] wire_363_1;
  assign wire_363 = wire_363_0|wire_363_1;
  wire [0:0] wire_364;
  wire [0:0] wire_365;
  wire [7:0] wire_366;
  wire [0:0] wire_367;
  wire [0:0] wire_368;
  wire [7:0] wire_369;
  wire [7:0] wire_370;
  wire [7:0] wire_371;
  wire [7:0] wire_372;
  wire [0:0] wire_373;
  wire [0:0] wire_374;
  wire [7:0] wire_375;
  wire [0:0] wire_376;
  wire [0:0] wire_377;
  wire [0:0] wire_378;
  wire [0:0] wire_379;
  wire [0:0] wire_380;
  wire [0:0] wire_381;
  wire [7:0] wire_382;
  wire [0:0] wire_383;
  wire [0:0] wire_384;
  wire [0:0] wire_385;
  wire [7:0] wire_386;
  wire [0:0] wire_387;
  wire [0:0] wire_388;
  wire [7:0] wire_389;
  wire [7:0] wire_390;
  wire [0:0] wire_391;
  wire [0:0] wire_392;
  wire [7:0] wire_393;
  wire [7:0] wire_394;
  wire [0:0] wire_395;
  wire [0:0] wire_396;
  wire [0:0] wire_397;
  wire [0:0] wire_398;
  wire [0:0] wire_399;
  wire [0:0] wire_400;
  wire [7:0] wire_401;
  wire [0:0] wire_402;
  wire [0:0] wire_403;
  wire [0:0] wire_404;
  wire [0:0] wire_405;
  wire [7:0] wire_406;
  wire [0:0] wire_407;
  wire [7:0] wire_408;
  wire [7:0] wire_409;
  wire [7:0] wire_410;
  wire [0:0] wire_411;
  wire [7:0] wire_412;
  wire [0:0] wire_413;
  wire [0:0] wire_414;
  wire [0:0] wire_415;
  wire [0:0] wire_416;
  wire [0:0] wire_417;
  wire [7:0] wire_418;
  wire [0:0] wire_419;
  wire [7:0] wire_420;
  wire [31:0] wire_421;
  wire [0:0] wire_422;
  wire [7:0] wire_423;
  wire [7:0] wire_424;
  wire [0:0] wire_425;
  wire [0:0] wire_426;
  wire [0:0] wire_427;
  wire [7:0] wire_428;
  wire [7:0] wire_429;
  wire [7:0] wire_430;
  wire [0:0] wire_431;
  wire [0:0] wire_432;
  wire [0:0] wire_433;
  wire [0:0] wire_434;
  wire [0:0] wire_435;
  wire [0:0] wire_436;
  wire [0:0] wire_437;
  wire [7:0] wire_438;

endmodule
