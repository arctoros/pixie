module Pixiez_Final (clk, rst, arch_output_enable, arch_output_value, arch_input_enable, arch_input_value);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;

  output  wire [0:0] arch_output_enable;
  output  wire [7:0] arch_output_value;
  output  wire [0:0] arch_input_enable;
  input  wire [7:0] arch_input_value;

  TC_Not # (.UUID(64'd680444558656414018 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_10), .out(wire_192));
  TC_Or3 # (.UUID(64'd534734424402985405 ^ UUID), .BIT_WIDTH(64'd1)) Or3_1 (.in0(wire_155), .in1(wire_176), .in2(wire_172), .out(wire_130));
  TC_Or3 # (.UUID(64'd4567130074526553310 ^ UUID), .BIT_WIDTH(64'd1)) Or3_2 (.in0(wire_174), .in1(wire_159), .in2(wire_58), .out(wire_212));
  TC_Or3 # (.UUID(64'd2737475285567390637 ^ UUID), .BIT_WIDTH(64'd1)) Or3_3 (.in0(wire_34), .in1(wire_118), .in2(wire_151), .out(wire_37));
  TC_Or3 # (.UUID(64'd1460121507051805330 ^ UUID), .BIT_WIDTH(64'd1)) Or3_4 (.in0(wire_37), .in1(wire_212), .in2(wire_205), .out(wire_144));
  TC_Not # (.UUID(64'd3263495404627770251 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_210), .out(wire_96));
  TC_DelayLine # (.UUID(64'd1861931133330004945 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_6 (.clk(clk), .rst(rst), .in(wire_96), .out(wire_210));
  TC_Not # (.UUID(64'd774824456586639901 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_161), .out(wire_97));
  TC_Or3 # (.UUID(64'd957665538453266802 ^ UUID), .BIT_WIDTH(64'd1)) Or3_8 (.in0(wire_112), .in1(wire_130), .in2(wire_169), .out(wire_161));
  TC_Add # (.UUID(64'd3301328818535174719 ^ UUID), .BIT_WIDTH(64'd8)) Add8_9 (.in0(wire_121), .in1(wire_133), .ci(wire_97), .out(wire_16), .co());
  TC_Or # (.UUID(64'd3186172645923730952 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_284), .in1(wire_291), .out(wire_155));
  TC_Not # (.UUID(64'd4418713765798495162 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_156), .out(wire_137));
  TC_Or3 # (.UUID(64'd3359031826937924206 ^ UUID), .BIT_WIDTH(64'd1)) Or3_12 (.in0(wire_4), .in1(wire_134), .in2(wire_231), .out(wire_284));
  TC_Decoder3 # (.UUID(64'd4465221940936740645 ^ UUID)) Decoder3_13 (.dis(wire_61), .sel0(wire_38[0:0]), .sel1(wire_164[0:0]), .sel2(wire_20[0:0]), .out0(wire_174), .out1(wire_152), .out2(wire_43), .out3(wire_234), .out4(wire_110), .out5(wire_89), .out6(wire_231), .out7(wire_160));
  TC_Decoder3 # (.UUID(64'd664854618839101163 ^ UUID)) Decoder3_14 (.dis(wire_256), .sel0(wire_38[0:0]), .sel1(wire_164[0:0]), .sel2(wire_20[0:0]), .out0(wire_28), .out1(wire_58), .out2(wire_159), .out3(wire_208), .out4(wire_298), .out5(wire_146), .out6(wire_50), .out7(wire_225));
  TC_Decoder3 # (.UUID(64'd388458847481545701 ^ UUID)) Decoder3_15 (.dis(wire_120), .sel0(wire_38[0:0]), .sel1(wire_164[0:0]), .sel2(wire_20[0:0]), .out0(wire_139), .out1(wire_9), .out2(wire_88), .out3(wire_65), .out4(wire_239), .out5(wire_51), .out6(wire_100), .out7(wire_17));
  TC_Decoder3 # (.UUID(64'd1325274093033025990 ^ UUID)) Decoder3_16 (.dis(wire_294), .sel0(wire_38[0:0]), .sel1(wire_164[0:0]), .sel2(wire_20[0:0]), .out0(wire_168), .out1(wire_151), .out2(wire_118), .out3(wire_34), .out4(wire_116), .out5(wire_268), .out6(wire_113), .out7(wire_18));
  TC_Not # (.UUID(64'd56215910927289989 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_173), .out(wire_61));
  TC_Not # (.UUID(64'd1568445558185814797 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_131), .out(wire_294));
  TC_Not # (.UUID(64'd3688819333690076749 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_232), .out(wire_120));
  TC_Not # (.UUID(64'd2914649659429896514 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_304), .out(wire_256));
  TC_Maker8 # (.UUID(64'd4274226248529413390 ^ UUID)) Maker8_21 (.in0(wire_174), .in1(wire_152), .in2(wire_43), .in3(wire_234), .in4(wire_110), .in5(wire_89), .in6(wire_231), .in7(wire_160), .out(wire_222));
  TC_Maker8 # (.UUID(64'd2503620967526902392 ^ UUID)) Maker8_22 (.in0(wire_28), .in1(wire_58), .in2(wire_159), .in3(wire_208), .in4(wire_298), .in5(wire_146), .in6(wire_50), .in7(wire_225), .out(wire_207));
  TC_Maker8 # (.UUID(64'd736697256551715288 ^ UUID)) Maker8_23 (.in0(wire_139), .in1(wire_9), .in2(wire_88), .in3(wire_65), .in4(wire_239), .in5(wire_51), .in6(wire_100), .in7(wire_17), .out(wire_274));
  TC_Maker8 # (.UUID(64'd832968618284013991 ^ UUID)) Maker8_24 (.in0(wire_168), .in1(wire_151), .in2(wire_118), .in3(wire_34), .in4(wire_116), .in5(wire_268), .in6(wire_113), .in7(wire_18), .out(wire_229));
  TC_Or3 # (.UUID(64'd2334335797361251671 ^ UUID), .BIT_WIDTH(64'd1)) Or3_25 (.in0(wire_50), .in1(wire_225), .in2(wire_234), .out(wire_134));
  TC_Or3 # (.UUID(64'd4505646521355499044 ^ UUID), .BIT_WIDTH(64'd1)) Or3_26 (.in0(wire_268), .in1(wire_18), .in2(wire_139), .out(wire_291));
  TC_Or3 # (.UUID(64'd2771484508194729184 ^ UUID), .BIT_WIDTH(64'd1)) Or3_27 (.in0(wire_51), .in1(wire_239), .in2(wire_65), .out(wire_283));
  TC_Or3 # (.UUID(64'd2848731522163985212 ^ UUID), .BIT_WIDTH(64'd1)) Or3_28 (.in0(wire_28), .in1(wire_17), .in2(wire_100), .out(wire_106));
  TC_DelayLine # (.UUID(64'd1068115119822942229 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_29 (.clk(clk), .rst(rst), .in(wire_11[7:0]), .out(wire_277));
  TC_DelayLine # (.UUID(64'd804044612046236745 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_227), .out(wire_10));
  TC_Splitter16 # (.UUID(64'd1875228578544666958 ^ UUID)) Splitter16_31 (.in(wire_238), .out0(wire_300), .out1(wire_25));
  TC_Maker16 # (.UUID(64'd3608744494562313405 ^ UUID)) Maker16_32 (.in0({{7{1'b0}}, wire_192 }), .in1(wire_189), .out(wire_238));
  TC_Or3 # (.UUID(64'd3746619389515595809 ^ UUID), .BIT_WIDTH(64'd1)) Or3_33 (.in0(wire_27), .in1(wire_29), .in2(wire_140), .out(wire_227));
  TC_Not # (.UUID(64'd966737772035534885 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_75[0:0]), .out(wire_228));
  TC_Not # (.UUID(64'd424140961992658426 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_57[0:0]), .out(wire_166));
  TC_Splitter32 # (.UUID(64'd2809680451032690949 ^ UUID)) Splitter32_36 (.in(wire_62), .out0(wire_290), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd2117984546099265654 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_37 (.out(wire_22));
  TC_Mux # (.UUID(64'd2353982102422779838 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_63), .in0(wire_5), .in1(wire_22), .out(wire_276));
  TC_Add # (.UUID(64'd4134817076244850895 ^ UUID), .BIT_WIDTH(64'd8)) Add8_39 (.in0(wire_6), .in1(wire_276), .ci(1'd0), .out(wire_204), .co());
  TC_Constant # (.UUID(64'd1952156418708934468 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_40 (.out(wire_191));
  TC_Mux # (.UUID(64'd4094225513381061300 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_41 (.sel(wire_66), .in0(wire_5), .in1(wire_191), .out(wire_301));
  TC_Neg # (.UUID(64'd102576365000716770 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_42 (.in(wire_301), .out(wire_285));
  TC_Add # (.UUID(64'd2689942381287690498 ^ UUID), .BIT_WIDTH(64'd8)) Add8_43 (.in0(wire_6), .in1(wire_285), .ci(1'd0), .out(wire_271), .co());
  TC_Switch # (.UUID(64'd4137287338459891824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_44 (.en(wire_254), .in(wire_271), .out(wire_11_8[7:0]));
  TC_Switch # (.UUID(64'd1351346083360514605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_105), .in(wire_204), .out(wire_11_11[7:0]));
  TC_Splitter8 # (.UUID(64'd4357406098891943912 ^ UUID)) Splitter8_46 (.in(wire_290), .out0(wire_206), .out1(wire_243), .out2(), .out3(), .out4(wire_48), .out5(wire_63), .out6(wire_66), .out7(wire_270));
  TC_Not # (.UUID(64'd3532098913873322011 ^ UUID), .BIT_WIDTH(64'd1)) Not_47 (.in(wire_71[0:0]), .out(wire_286));
  TC_Switch # (.UUID(64'd2937048381182156076 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_48 (.en(wire_156), .in(wire_95), .out(wire_6_18));
  TC_Switch # (.UUID(64'd412107824868226985 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_49 (.en(wire_137), .in(wire_95), .out(wire_145));
  TC_Switch # (.UUID(64'd1458121506772114657 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_75[0:0]), .in(wire_72), .out(wire_5_1));
  TC_Switch # (.UUID(64'd2507210810598866832 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_228), .in(wire_72), .out(wire_175));
  TC_Switch # (.UUID(64'd1855204595012977435 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_71[0:0]), .in(wire_91), .out(wire_11_5[7:0]));
  TC_Switch # (.UUID(64'd1879885438156656135 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_286), .in(wire_91), .out(wire_13));
  TC_Splitter16 # (.UUID(64'd4592662178931061204 ^ UUID)) Splitter16_54 (.in(wire_224), .out0(wire_44), .out1(wire_57));
  TC_Or3 # (.UUID(64'd1577578265915915529 ^ UUID), .BIT_WIDTH(64'd1)) Or3_55 (.in0(wire_44[0:0]), .in1(wire_57[0:0]), .in2(wire_112), .out(wire_132));
  TC_Switch # (.UUID(64'd2610614871112416436 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_56 (.en(wire_44[0:0]), .in(wire_54[7:0]), .out(wire_299));
  TC_Switch # (.UUID(64'd165300680693317419 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_57 (.en(wire_44[0:0]), .in(wire_261[7:0]), .out(wire_72));
  TC_Switch # (.UUID(64'd2260740780324363689 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_58 (.en(wire_132), .in(wire_297[7:0]), .out(wire_95));
  TC_Mux # (.UUID(64'd4528590367296190010 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_59 (.sel(wire_166), .in0(wire_261[7:0]), .in1(wire_299), .out(wire_91));
  TC_Splitter16 # (.UUID(64'd2701914707745210702 ^ UUID)) Splitter16_60 (.in(wire_278), .out0(wire_71), .out1(wire_75));
  TC_Maker16 # (.UUID(64'd1365218859602849489 ^ UUID)) Maker16_61 (.in0({{7{1'b0}}, wire_255 }), .in1({{7{1'b0}}, wire_272 }), .out(wire_278));
  TC_Switch # (.UUID(64'd2155635750972134594 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_62 (.en(wire_10), .in(wire_277), .out(wire_189));
  TC_Mux # (.UUID(64'd1791751815309933921 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_63 (.sel(wire_300[0:0]), .in0(wire_25), .in1(wire_198), .out(wire_121));
  TC_Maker16 # (.UUID(64'd3395313277560932739 ^ UUID)) Maker16_64 (.in0({{7{1'b0}}, wire_169 }), .in1({{7{1'b0}}, wire_130 }), .out(wire_224));
  TC_Not # (.UUID(64'd3453103485371531751 ^ UUID), .BIT_WIDTH(64'd1)) Not_65 (.in(wire_96), .out(wire_233));
  TC_Counter # (.UUID(64'd1171561396707692790 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_66 (.clk(clk), .rst(rst), .save(wire_96), .in(wire_16), .out(wire_248));
  TC_Counter # (.UUID(64'd2621291279726673638 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_67 (.clk(clk), .rst(rst), .save(wire_210), .in(wire_16), .out(wire_279));
  TC_Switch # (.UUID(64'd1839974249620431880 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_68 (.en(wire_233), .in(wire_248), .out(wire_198_0));
  TC_Switch # (.UUID(64'd1170108399670313272 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_69 (.en(wire_96), .in(wire_279), .out(wire_198_1));
  TC_Constant # (.UUID(64'd358007510611002277 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_70 (.out(wire_260));
  TC_Constant # (.UUID(64'd3874548421935569254 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_71 (.out(wire_218));
  TC_Constant # (.UUID(64'd1203375723678859801 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_72 (.out(wire_306));
  TC_Switch # (.UUID(64'd1933124139798812111 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_73 (.en(wire_112), .in(wire_260), .out(wire_133_2));
  TC_Switch # (.UUID(64'd287643768980040071 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_74 (.en(wire_130), .in(wire_218), .out(wire_133_0));
  TC_Switch # (.UUID(64'd4195386940103341620 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_169), .in(wire_306), .out(wire_133_1));
  TC_Splitter8 # (.UUID(64'd2599557092287595297 ^ UUID)) Splitter8_76 (.in(wire_165[7:0]), .out0(wire_293), .out1(wire_308), .out2(wire_80), .out3(wire_259), .out4(wire_264), .out5(wire_255), .out6(wire_272), .out7(wire_156));
  TC_Ram # (.UUID(64'd1708105537810654235 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_77 (.clk(clk), .rst(rst), .load(wire_196), .save(wire_1), .address({{24{1'b0}}, wire_5 }), .in0({{56{1'b0}}, wire_6 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_11_2), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd97660009947370162 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd128)) Ram_78 (.clk(clk), .rst(rst), .load(wire_47), .save(wire_68), .address({{24{1'b0}}, wire_85 }), .in0({{56{1'b0}}, wire_16 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_281), .out1(), .out2(), .out3());
  TC_Or # (.UUID(64'd733084299857471502 ^ UUID), .BIT_WIDTH(64'd1)) Or_79 (.in0(wire_68), .in1(wire_47), .out(wire_29));
  TC_Splitter32 # (.UUID(64'd3048987527585864498 ^ UUID)) Splitter32_80 (.in(wire_62), .out0(), .out1(wire_40), .out2(), .out3(wire_41));
  TC_Or # (.UUID(64'd4064324485441264957 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_47), .in1(wire_68), .out(wire_125));
  TC_Switch # (.UUID(64'd2955305895674404779 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_82 (.en(wire_47), .in(wire_281[7:0]), .out(wire_11_7[7:0]));
  TC_Switch # (.UUID(64'd3592902196704226444 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_83 (.en(wire_68), .in(wire_6), .out(wire_11_4[7:0]));
  TC_Register # (.UUID(64'd4471884361578131577 ^ UUID), .BIT_WIDTH(64'd8)) Register8_84 (.clk(clk), .rst(rst), .load(wire_125), .save(wire_125), .in(wire_214), .out(wire_84));
  TC_Switch # (.UUID(64'd4562232227874677430 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_85 (.en(wire_68), .in(wire_30), .out(wire_214_0));
  TC_Switch # (.UUID(64'd114510401986147547 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_86 (.en(wire_68), .in(wire_214), .out(wire_85_0));
  TC_Add # (.UUID(64'd263770477141513169 ^ UUID), .BIT_WIDTH(64'd8)) Add8_87 (.in0(wire_81), .in1(wire_84), .ci(1'd0), .out(wire_30), .co());
  TC_Switch # (.UUID(64'd2865125256828769888 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_88 (.en(wire_47), .in(wire_302), .out(wire_214_1));
  TC_Switch # (.UUID(64'd1945149825988830027 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_89 (.en(wire_47), .in(wire_84), .out(wire_85_1));
  TC_Constant # (.UUID(64'd2864754851009931669 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_90 (.out(wire_81));
  TC_Neg # (.UUID(64'd1766191137768834313 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_91 (.in(wire_81), .out(wire_250));
  TC_Add # (.UUID(64'd1197352873015043648 ^ UUID), .BIT_WIDTH(64'd8)) Add8_92 (.in0(wire_84), .in1(wire_250), .ci(1'd0), .out(wire_302), .co());
  TC_Splitter8 # (.UUID(64'd3473615707126412287 ^ UUID)) Splitter8_93 (.in(wire_41), .out0(wire_1), .out1(wire_196), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_46));
  TC_Constant # (.UUID(64'd3007591360524826255 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_94 (.out(wire_163));
  TC_Or # (.UUID(64'd3353986015329929110 ^ UUID), .BIT_WIDTH(64'd1)) Or_95 (.in0(wire_128), .in1(wire_142), .out(wire_295));
  TC_LessU # (.UUID(64'd2857803572762207218 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_96 (.in0(wire_5), .in1(wire_6), .out(wire_142));
  TC_Not # (.UUID(64'd3713135576456282771 ^ UUID), .BIT_WIDTH(64'd1)) Not_97 (.in(wire_128), .out(wire_230));
  TC_Or # (.UUID(64'd1283831029887634373 ^ UUID), .BIT_WIDTH(64'd1)) Or_98 (.in0(wire_111), .in1(wire_128), .out(wire_53));
  TC_Equal # (.UUID(64'd3249866343864622854 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_99 (.in0(wire_6), .in1(wire_5), .out(wire_128));
  TC_LessU # (.UUID(64'd2949327424893302673 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_100 (.in0(wire_6), .in1(wire_5), .out(wire_111));
  TC_Equal # (.UUID(64'd3467215832225421993 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_101 (.in0(wire_163), .in1(wire_6), .out(wire_267));
  TC_Constant # (.UUID(64'd4251321236624205294 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_102 (.out(wire_220));
  TC_Switch # (.UUID(64'd4268044874154730043 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_103 (.en(wire_226), .in(wire_220), .out(wire_140_5));
  TC_Switch # (.UUID(64'd1386783397630713083 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_104 (.en(wire_138), .in(wire_267), .out(wire_140_3));
  TC_Switch # (.UUID(64'd1155028069485320511 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_105 (.en(wire_251), .in(wire_111), .out(wire_140_0));
  TC_Switch # (.UUID(64'd3348470806054818924 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_106 (.en(wire_199), .in(wire_53), .out(wire_140_1));
  TC_Switch # (.UUID(64'd1041869814803847902 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_107 (.en(wire_24), .in(wire_128), .out(wire_140_2));
  TC_Switch # (.UUID(64'd4055918702281020749 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_108 (.en(wire_245), .in(wire_230), .out(wire_140_4));
  TC_Switch # (.UUID(64'd3083535767069260986 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_109 (.en(wire_237), .in(wire_295), .out(wire_140_6));
  TC_Switch # (.UUID(64'd2913504031160566908 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_110 (.en(wire_242), .in(wire_142), .out(wire_140_7));
  TC_Splitter8 # (.UUID(64'd1194059391229914692 ^ UUID)) Splitter8_111 (.in(wire_40), .out0(wire_226), .out1(wire_138), .out2(wire_251), .out3(wire_199), .out4(wire_24), .out5(wire_245), .out6(wire_237), .out7(wire_242));
  TC_Register # (.UUID(64'd1786549938381629068 ^ UUID), .BIT_WIDTH(64'd8)) Register8_112 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_188), .in(wire_11[7:0]), .out(wire_56));
  TC_Register # (.UUID(64'd2601905860340903537 ^ UUID), .BIT_WIDTH(64'd8)) Register8_113 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_190), .in(wire_11[7:0]), .out(wire_180));
  TC_Register # (.UUID(64'd2818150811460271121 ^ UUID), .BIT_WIDTH(64'd8)) Register8_114 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_23), .in(wire_11[7:0]), .out(wire_183));
  TC_Register # (.UUID(64'd3810474016475870525 ^ UUID), .BIT_WIDTH(64'd8)) Register8_115 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_167), .in(wire_11[7:0]), .out(wire_201));
  TC_Register # (.UUID(64'd1636002980180907684 ^ UUID), .BIT_WIDTH(64'd8)) Register8_116 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_249), .in(wire_11[7:0]), .out(wire_269));
  TC_Register # (.UUID(64'd3256658416273011892 ^ UUID), .BIT_WIDTH(64'd8)) Register8_117 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_141), .in(wire_11[7:0]), .out(wire_73));
  TC_Register # (.UUID(64'd2526494128293687363 ^ UUID), .BIT_WIDTH(64'd8)) Register8_118 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_83), .in(wire_11[7:0]), .out(wire_177));
  TC_Register # (.UUID(64'd3472073544120575095 ^ UUID), .BIT_WIDTH(64'd8)) Register8_119 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_76), .in(wire_11[7:0]), .out(wire_171));
  TC_Register # (.UUID(64'd542285582491664182 ^ UUID), .BIT_WIDTH(64'd8)) Register8_120 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_98), .in(wire_11[7:0]), .out(wire_148));
  TC_Register # (.UUID(64'd2124618488310653916 ^ UUID), .BIT_WIDTH(64'd8)) Register8_121 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_178), .in(wire_11[7:0]), .out(wire_49));
  TC_Register # (.UUID(64'd240222191994770064 ^ UUID), .BIT_WIDTH(64'd8)) Register8_122 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_122), .in(wire_11[7:0]), .out(wire_158));
  TC_Switch # (.UUID(64'd2919893529833212573 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_123 (.en(wire_129), .in(wire_183), .out(wire_6_17));
  TC_Switch # (.UUID(64'd2892052628952263194 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_124 (.en(wire_236), .in(wire_183), .out(wire_32_11));
  TC_Switch # (.UUID(64'd1045466942081498185 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_125 (.en(wire_257), .in(wire_201), .out(wire_6_16));
  TC_Switch # (.UUID(64'd4352568465751771503 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_126 (.en(wire_162), .in(wire_201), .out(wire_32_9));
  TC_Switch # (.UUID(64'd294837876173931186 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_127 (.en(wire_103), .in(wire_177), .out(wire_6_15));
  TC_Switch # (.UUID(64'd718804107324007425 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_128 (.en(wire_149), .in(wire_177), .out(wire_32_7));
  TC_Switch # (.UUID(64'd2106337721725300490 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_129 (.en(wire_8), .in(wire_148), .out(wire_6_13));
  TC_Switch # (.UUID(64'd1382626067278158580 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_130 (.en(wire_153), .in(wire_148), .out(wire_32_5));
  TC_Switch # (.UUID(64'd4280389427710179554 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_131 (.en(wire_240), .in(wire_171), .out(wire_6_12));
  TC_Switch # (.UUID(64'd2870197787210989981 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_132 (.en(wire_86), .in(wire_171), .out(wire_32_3));
  TC_Switch # (.UUID(64'd1025076596807518358 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_133 (.en(wire_31), .in(wire_269), .out(wire_6_10));
  TC_Switch # (.UUID(64'd961920732700576390 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_134 (.en(wire_266), .in(wire_269), .out(wire_32_1));
  TC_Switch # (.UUID(64'd455633754159767112 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_135 (.en(wire_262), .in(wire_49), .out(wire_6_8));
  TC_Switch # (.UUID(64'd3572372897415253218 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_136 (.en(wire_87), .in(wire_49), .out(wire_32_0));
  TC_Switch # (.UUID(64'd2693638907193452534 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_137 (.en(wire_135), .in(wire_73), .out(wire_6_6));
  TC_Switch # (.UUID(64'd4344217990313000347 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_138 (.en(wire_19), .in(wire_73), .out(wire_32_2));
  TC_Switch # (.UUID(64'd258289412669476303 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_139 (.en(wire_104), .in(wire_180), .out(wire_6_4));
  TC_Switch # (.UUID(64'd4506884556720173301 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_140 (.en(wire_12), .in(wire_180), .out(wire_32_4));
  TC_Switch # (.UUID(64'd3160999002775359256 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_141 (.en(wire_235), .in(wire_56), .out(wire_6_2));
  TC_Switch # (.UUID(64'd4258632307214665985 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_142 (.en(wire_93), .in(wire_56), .out(wire_32_6));
  TC_Switch # (.UUID(64'd1115547685276398812 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_143 (.en(wire_197), .in(wire_158), .out(wire_6_0));
  TC_Switch # (.UUID(64'd2594916914153554215 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_144 (.en(wire_82), .in(wire_158), .out(wire_32_8));
  TC_Switch # (.UUID(64'd2067768058777429209 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_145 (.en(wire_7), .in(wire_74), .out(wire_32_12));
  TC_Switch # (.UUID(64'd1049797112137663963 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_146 (.en(wire_193), .in(wire_74), .out(wire_6_3));
  TC_Switch # (.UUID(64'd4067917907888700042 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_147 (.en(wire_247), .in(wire_67), .out(wire_32_10));
  TC_Switch # (.UUID(64'd3311537942366866912 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_148 (.en(wire_33), .in(wire_67), .out(wire_6_1));
  TC_Register # (.UUID(64'd1377807017811864986 ^ UUID), .BIT_WIDTH(64'd8)) Register8_149 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_195), .in(wire_11[7:0]), .out(wire_67));
  TC_Register # (.UUID(64'd1236368519178447850 ^ UUID), .BIT_WIDTH(64'd8)) Register8_150 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_157), .in(wire_11[7:0]), .out(wire_74));
  TC_Splitter8 # (.UUID(64'd2271575679199078636 ^ UUID)) Splitter8_151 (.in(wire_127), .out0(), .out1(), .out2(wire_14), .out3(wire_45), .out4(wire_68), .out5(wire_47), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd261396410293330702 ^ UUID)) Splitter32_152 (.in(wire_62), .out0(), .out1(), .out2(), .out3(wire_127));
  TC_Ram # (.UUID(64'd4117401978527469154 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd32)) Ram_153 (.clk(clk), .rst(rst), .load(wire_45), .save(wire_14), .address({{24{1'b0}}, wire_221 }), .in0({{56{1'b0}}, wire_6 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_11_0), .out1(), .out2(), .out3());
  TC_Switch # (.UUID(64'd3161290829479641019 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_154 (.en(wire_48), .in(wire_102), .out(wire_11_6[7:0]));
  TC_Switch # (.UUID(64'd3115314308242652354 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_155 (.en(wire_270), .in(wire_217), .out(wire_11_3[7:0]));
  TC_Neg # (.UUID(64'd77226668367061539 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_156 (.in(wire_6), .out(wire_102));
  TC_Or # (.UUID(64'd1380170131908116772 ^ UUID), .BIT_WIDTH(64'd1)) Or_157 (.in0(wire_66), .in1(wire_243), .out(wire_254));
  TC_Constant # (.UUID(64'd1678158762324492118 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_158 (.out(wire_64));
  TC_Ashr # (.UUID(64'd1558764338386234982 ^ UUID), .BIT_WIDTH(64'd8)) Ashr8_159 (.in(wire_6), .shift(wire_64), .out(wire_217));
  TC_Constant # (.UUID(64'd2997253212554120558 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_160 (.out(wire_2));
  TC_Constant # (.UUID(64'd3797620182831446698 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_161 (.out(wire_252));
  TC_Neg # (.UUID(64'd3558537661740369771 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_162 (.in(wire_252), .out(wire_307));
  TC_Register # (.UUID(64'd2759537605007938592 ^ UUID), .BIT_WIDTH(64'd8)) Register8_163 (.clk(clk), .rst(rst), .load(wire_170), .save(wire_170), .in(wire_184), .out(wire_69));
  TC_Switch # (.UUID(64'd929829793202303828 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_164 (.en(wire_14), .in(wire_187), .out(wire_184_1));
  TC_Switch # (.UUID(64'd3728124673178845213 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_165 (.en(wire_14), .in(wire_184), .out(wire_221_1));
  TC_Add # (.UUID(64'd1902099203606853874 ^ UUID), .BIT_WIDTH(64'd8)) Add8_166 (.in0(wire_252), .in1(wire_69), .ci(1'd0), .out(wire_187), .co());
  TC_Switch # (.UUID(64'd3498208789273416986 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_167 (.en(wire_45), .in(wire_109), .out(wire_184_0));
  TC_Switch # (.UUID(64'd1321154288873073244 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_168 (.en(wire_45), .in(wire_69), .out(wire_221_0));
  TC_Or # (.UUID(64'd1321825518205599775 ^ UUID), .BIT_WIDTH(64'd1)) Or_169 (.in0(wire_45), .in1(wire_14), .out(wire_170));
  TC_Add # (.UUID(64'd4199771119303044950 ^ UUID), .BIT_WIDTH(64'd8)) Add8_170 (.in0(wire_69), .in1(wire_307), .ci(1'd0), .out(wire_109), .co());
  TC_Switch # (.UUID(64'd81193405753331740 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_171 (.en(wire_186), .in(wire_273), .out(wire_11_17[7:0]));
  TC_Switch # (.UUID(64'd4415608983622849585 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_172 (.en(wire_202), .in(wire_115), .out(wire_11_16[7:0]));
  TC_And # (.UUID(64'd1669263777784106749 ^ UUID), .BIT_WIDTH(64'd8)) And8_173 (.in0(wire_6), .in1(wire_5), .out(wire_273));
  TC_Or # (.UUID(64'd873622160744398625 ^ UUID), .BIT_WIDTH(64'd8)) Or8_174 (.in0(wire_6), .in1(wire_5), .out(wire_115));
  TC_Xor # (.UUID(64'd2690694932656199993 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_175 (.in0(wire_6), .in1(wire_5), .out(wire_123));
  TC_Not # (.UUID(64'd3218967706620565239 ^ UUID), .BIT_WIDTH(64'd8)) Not8_176 (.in(wire_6), .out(wire_154));
  TC_Shl # (.UUID(64'd3160996752802486419 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_177 (.in(wire_6), .shift({{7{1'b0}}, wire_108 }), .out(wire_280));
  TC_Shr # (.UUID(64'd1938059414175291844 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_178 (.in(wire_6), .shift({{7{1'b0}}, wire_108 }), .out(wire_296));
  TC_Rol # (.UUID(64'd379560068498716864 ^ UUID), .BIT_WIDTH(64'd8)) Rol8_179 (.in(wire_6), .shift({{7{1'b0}}, wire_108 }), .out(wire_244));
  TC_Ror # (.UUID(64'd4299448326393726552 ^ UUID), .BIT_WIDTH(64'd8)) Ror8_180 (.in(wire_6), .shift({{7{1'b0}}, wire_108 }), .out(wire_194));
  TC_Switch # (.UUID(64'd2309803132069263134 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_181 (.en(wire_182), .in(wire_123), .out(wire_11_15[7:0]));
  TC_Switch # (.UUID(64'd2923996340214116429 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_182 (.en(wire_263), .in(wire_154), .out(wire_11_14[7:0]));
  TC_Switch # (.UUID(64'd2407013580594625997 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_183 (.en(wire_36), .in(wire_296), .out(wire_11_13[7:0]));
  TC_Switch # (.UUID(64'd3621734594009664278 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_184 (.en(wire_126), .in(wire_280), .out(wire_11_12[7:0]));
  TC_Switch # (.UUID(64'd1878036650580289106 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_185 (.en(wire_213), .in(wire_194), .out(wire_11_10[7:0]));
  TC_Switch # (.UUID(64'd4077902765271428258 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_186 (.en(wire_282), .in(wire_244), .out(wire_11_9[7:0]));
  TC_Splitter8 # (.UUID(64'd772965213957027290 ^ UUID)) Splitter8_187 (.in(wire_216), .out0(wire_186), .out1(wire_202), .out2(wire_182), .out3(wire_263), .out4(wire_36), .out5(wire_126), .out6(wire_213), .out7(wire_282));
  TC_Splitter32 # (.UUID(64'd3454244281776476436 ^ UUID)) Splitter32_188 (.in(wire_62), .out0(), .out1(), .out2(wire_216), .out3());
  TC_Register # (.UUID(64'd1044465739269958273 ^ UUID), .BIT_WIDTH(64'd8)) Register8_189 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_52), .in(wire_11[7:0]), .out(wire_143));
  TC_Register # (.UUID(64'd1014775350705063680 ^ UUID), .BIT_WIDTH(64'd8)) Register8_190 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_150), .in(wire_11[7:0]), .out(wire_117));
  TC_Switch # (.UUID(64'd17400449972985902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_191 (.en(wire_92), .in(wire_117), .out(wire_6_5));
  TC_Switch # (.UUID(64'd1757317349619379473 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_192 (.en(wire_211), .in(wire_117), .out(wire_32_13));
  TC_Switch # (.UUID(64'd347935731390232235 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_193 (.en(wire_287), .in(wire_143), .out(wire_6_7));
  TC_Switch # (.UUID(64'd347572746678109137 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_194 (.en(wire_101), .in(wire_143), .out(wire_32_14));
  TC_Not # (.UUID(64'd2075639373923651350 ^ UUID), .BIT_WIDTH(64'd1)) Not_195 (.in(wire_78), .out(wire_0));
  TC_And # (.UUID(64'd754894496948066040 ^ UUID), .BIT_WIDTH(64'd1)) And_196 (.in0(wire_78), .in1(wire_42), .out(wire_241));
  TC_Or # (.UUID(64'd805549193662201184 ^ UUID), .BIT_WIDTH(64'd1)) Or_197 (.in0(wire_42), .in1(wire_0), .out(wire_99));
  TC_Decoder3 # (.UUID(64'd3761069498695685674 ^ UUID)) Decoder3_198 (.dis(wire_136), .sel0(wire_59), .sel1(wire_94), .sel2(wire_185), .out0(wire_129), .out1(wire_257), .out2(wire_103), .out3(wire_8), .out4(wire_240), .out5(wire_31), .out6(wire_262), .out7(wire_135));
  TC_Decoder3 # (.UUID(64'd1604216519862450208 ^ UUID)) Decoder3_199 (.dis(wire_99), .sel0(wire_59), .sel1(wire_94), .sel2(wire_185), .out0(wire_104), .out1(wire_235), .out2(wire_197), .out3(wire_33), .out4(wire_193), .out5(wire_92), .out6(wire_287), .out7(wire_288));
  TC_Or # (.UUID(64'd259192617280007518 ^ UUID), .BIT_WIDTH(64'd1)) Or_200 (.in0(wire_26), .in1(wire_253), .out(wire_258));
  TC_Decoder3 # (.UUID(64'd1295781503081853777 ^ UUID)) Decoder3_201 (.dis(wire_77), .sel0(wire_35), .sel1(wire_70), .sel2(wire_21), .out0(wire_236), .out1(wire_162), .out2(wire_149), .out3(wire_153), .out4(wire_86), .out5(wire_266), .out6(wire_87), .out7(wire_19));
  TC_Decoder3 # (.UUID(64'd57268074239693712 ^ UUID)) Decoder3_202 (.dis(wire_258), .sel0(wire_35), .sel1(wire_70), .sel2(wire_21), .out0(wire_12), .out1(wire_93), .out2(wire_82), .out3(wire_247), .out4(wire_7), .out5(wire_211), .out6(wire_101), .out7(wire_223));
  TC_Or # (.UUID(64'd1404831056388826959 ^ UUID), .BIT_WIDTH(64'd1)) Or_203 (.in0(wire_3), .in1(wire_124), .out(wire_292));
  TC_And # (.UUID(64'd2552562799264486541 ^ UUID), .BIT_WIDTH(64'd1)) And_204 (.in0(wire_179), .in1(wire_3), .out(wire_107));
  TC_Decoder3 # (.UUID(64'd762150619108810778 ^ UUID)) Decoder3_205 (.dis(wire_292), .sel0(wire_275), .sel1(wire_119), .sel2(wire_15), .out0(wire_190), .out1(wire_188), .out2(wire_122), .out3(wire_195), .out4(wire_157), .out5(wire_150), .out6(wire_52), .out7(wire_181));
  TC_Decoder3 # (.UUID(64'd494457670381439667 ^ UUID)) Decoder3_206 (.dis(wire_60), .sel0(wire_275), .sel1(wire_119), .sel2(wire_15), .out0(wire_23), .out1(wire_167), .out2(wire_83), .out3(wire_98), .out4(wire_76), .out5(wire_249), .out6(wire_178), .out7(wire_141));
  TC_Splitter8 # (.UUID(64'd448586870420520821 ^ UUID)) Splitter8_207 (.in(wire_13), .out0(wire_275), .out1(wire_119), .out2(wire_15), .out3(wire_179), .out4(wire_3), .out5(), .out6(), .out7());
  TC_Or3 # (.UUID(64'd1235965720506732026 ^ UUID), .BIT_WIDTH(64'd1)) Or3_208 (.in0(wire_106), .in1(wire_283), .in2(wire_209), .out(wire_205));
  TC_Or3 # (.UUID(64'd64656781117703189 ^ UUID), .BIT_WIDTH(64'd1)) Or3_209 (.in0(wire_200[0:0]), .in1(wire_90), .in2(wire_26), .out(wire_77));
  TC_Not # (.UUID(64'd3756682246155706392 ^ UUID), .BIT_WIDTH(64'd1)) Not_210 (.in(wire_179), .out(wire_124));
  TC_Or3 # (.UUID(64'd1985979777212458751 ^ UUID), .BIT_WIDTH(64'd1)) Or3_211 (.in0(wire_289), .in1(wire_71[0:0]), .in2(wire_215), .out(wire_60));
  TC_Or3 # (.UUID(64'd1657864677517986892 ^ UUID), .BIT_WIDTH(64'd1)) Or3_212 (.in0(wire_246[0:0]), .in1(wire_78), .in2(wire_42), .out(wire_136));
  TC_And # (.UUID(64'd422870372255371239 ^ UUID), .BIT_WIDTH(64'd1)) And_213 (.in0(wire_124), .in1(wire_3), .out(wire_27));
  TC_Splitter8 # (.UUID(64'd760659632282220270 ^ UUID)) Splitter8_214 (.in(wire_175), .out0(wire_35), .out1(wire_70), .out2(wire_21), .out3(wire_90), .out4(wire_26), .out5(), .out6(), .out7());
  TC_Splitter8 # (.UUID(64'd638362282452151696 ^ UUID)) Splitter8_215 (.in(wire_145), .out0(wire_59), .out1(wire_94), .out2(wire_185), .out3(wire_78), .out4(wire_42), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd3337535575473260291 ^ UUID), .BIT_WIDTH(64'd1)) And_216 (.in0(wire_42), .in1(wire_305), .out(wire_147));
  TC_Not # (.UUID(64'd558454314996824891 ^ UUID), .BIT_WIDTH(64'd1)) Not_217 (.in(wire_78), .out(wire_305));
  TC_Maker32 # (.UUID(64'd1972774908657050676 ^ UUID)) Maker32_218 (.in0(wire_229), .in1(wire_274), .in2(wire_207), .in3(wire_222), .out(wire_62));
  TC_Or # (.UUID(64'd2498810294022311638 ^ UUID), .BIT_WIDTH(64'd1)) Or_219 (.in0(wire_63), .in1(wire_206), .out(wire_105));
  TC_Switch # (.UUID(64'd2854933611415915645 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_220 (.en(wire_46), .in(wire_6), .out(wire_11_1[7:0]));
  TC_Or3 # (.UUID(64'd4211290242648182257 ^ UUID), .BIT_WIDTH(64'd1)) Or3_221 (.in0(wire_43), .in1(wire_110), .in2(wire_89), .out(wire_112));
  TC_Or # (.UUID(64'd4406510584467674262 ^ UUID), .BIT_WIDTH(64'd1)) Or_222 (.in0(wire_110), .in1(wire_89), .out(wire_289));
  TC_Or # (.UUID(64'd240802604651373700 ^ UUID), .BIT_WIDTH(64'd1)) Or_223 (.in0(wire_179), .in1(wire_3), .out(wire_215));
  TC_And # (.UUID(64'd647954593887269646 ^ UUID), .BIT_WIDTH(64'd1)) And_224 (.in0(wire_90), .in1(wire_26), .out(wire_219));
  TC_Splitter16 # (.UUID(64'd2940418270800807678 ^ UUID)) Splitter16_225 (.in(wire_55), .out0(wire_200), .out1(wire_246));
  TC_Maker16 # (.UUID(64'd4473516211661289785 ^ UUID)) Maker16_226 (.in0(wire_75), .in1({{7{1'b0}}, wire_156 }), .out(wire_55));
  TC_Or3 # (.UUID(64'd1738768736642702813 ^ UUID), .BIT_WIDTH(64'd1)) Or3_227 (.in0(wire_208), .in1(wire_298), .in2(wire_146), .out(wire_4));
  TC_Program # (.UUID(64'd145079491480902460 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2036D0761E9DB3C.w8.bin"), .ARG_SIG("Program_2036D0761E9DB3C=%s")) Program_228 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_121 }), .out0(wire_165), .out1(wire_297), .out2(wire_261), .out3(wire_54));
  TC_Not # (.UUID(64'd2924370506823732469 ^ UUID), .BIT_WIDTH(64'd1)) Not_229 (.in(wire_90), .out(wire_253));
  TC_Maker32 # (.UUID(64'd3731905900420244009 ^ UUID)) Maker32_230 (.in0({{7{1'b0}}, wire_293 }), .in1({{7{1'b0}}, wire_308 }), .in2({{7{1'b0}}, wire_80 }), .in3({{7{1'b0}}, wire_259 }), .out(wire_203));
  TC_Splitter32 # (.UUID(64'd3952628877771949754 ^ UUID)) Splitter32_231 (.in(wire_203), .out0(wire_38), .out1(wire_164), .out2(wire_20), .out3(wire_114));
  TC_Or # (.UUID(64'd1464181653386223728 ^ UUID), .BIT_WIDTH(64'd1)) Or_232 (.in0(wire_113), .in1(wire_116), .out(wire_172));
  TC_Or # (.UUID(64'd1071650078955089329 ^ UUID), .BIT_WIDTH(64'd1)) Or_233 (.in0(wire_88), .in1(wire_168), .out(wire_209));
  TC_Or # (.UUID(64'd3984947405899213483 ^ UUID), .BIT_WIDTH(64'd1)) Or_234 (.in0(wire_152), .in1(wire_144), .out(wire_169));
  TC_Or # (.UUID(64'd19590702580144813 ^ UUID), .BIT_WIDTH(64'd1)) Or_235 (.in0(wire_9), .in1(wire_160), .out(wire_176));
  TC_Decoder2 # (.UUID(64'd2363697850107914081 ^ UUID)) Decoder2_236 (.sel0(wire_114[0:0]), .sel1(wire_264), .out0(wire_131), .out1(wire_232), .out2(wire_304), .out3(wire_173));
  TC_Switch # (.UUID(64'd1090992316792881700 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_237 (.en(wire_288), .in(wire_265), .out(wire_6_9));
  TC_Switch # (.UUID(64'd4578422426788892621 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_238 (.en(wire_223), .in(wire_265), .out(wire_5_3));
  TC_Switch # (.UUID(64'd2981244423840958363 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_239 (.en(wire_241), .in(wire_39), .out(wire_6_11));
  TC_Switch # (.UUID(64'd4233253593413734408 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_240 (.en(wire_219), .in(wire_39), .out(wire_5_2));
  TC_Switch # (.UUID(64'd323511192384597787 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_241 (.en(wire_147), .in(wire_16), .out(wire_6_14));
  TC_IOSwitch # (.UUID(64'd1626475142369920112 ^ UUID), .BIT_WIDTH(64'd8)) LevelOutputArch_242 (.in(wire_11[7:0]), .en(wire_107), .out(arch_output_value));
  TC_Switch # (.UUID(64'd3868416457659096598 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_243 (.en(wire_79), .in(wire_16), .out(wire_5_0));
  TC_Register # (.UUID(64'd799015932801999712 ^ UUID), .BIT_WIDTH(64'd8)) Register8_244 (.clk(clk), .rst(rst), .load(wire_2), .save(wire_181), .in(wire_11[7:0]), .out(wire_265));
  TC_Switch # (.UUID(64'd974745753494790983 ^ UUID), .BIT_WIDTH(64'd8)) LevelInputArch_245 (.en(wire_2), .in(arch_input_value), .out(wire_39));
  TC_And # (.UUID(64'd2334144837756105628 ^ UUID), .BIT_WIDTH(64'd1)) And_246 (.in0(wire_26), .in1(wire_303), .out(wire_79));
  TC_Not # (.UUID(64'd2110701898339003391 ^ UUID), .BIT_WIDTH(64'd1)) Not_247 (.in(wire_90), .out(wire_303));
  TC_Constant # (.UUID(64'd2996855662000809421 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_248 (.out(wire_108));

  wire [0:0] wire_0;
  wire [0:0] wire_1;
  wire [0:0] wire_2;
  assign arch_input_enable = wire_2;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [7:0] wire_5;
  wire [7:0] wire_5_0;
  wire [7:0] wire_5_1;
  wire [7:0] wire_5_2;
  wire [7:0] wire_5_3;
  assign wire_5 = wire_5_0|wire_5_1|wire_5_2|wire_5_3;
  wire [7:0] wire_6;
  wire [7:0] wire_6_0;
  wire [7:0] wire_6_1;
  wire [7:0] wire_6_2;
  wire [7:0] wire_6_3;
  wire [7:0] wire_6_4;
  wire [7:0] wire_6_5;
  wire [7:0] wire_6_6;
  wire [7:0] wire_6_7;
  wire [7:0] wire_6_8;
  wire [7:0] wire_6_9;
  wire [7:0] wire_6_10;
  wire [7:0] wire_6_11;
  wire [7:0] wire_6_12;
  wire [7:0] wire_6_13;
  wire [7:0] wire_6_14;
  wire [7:0] wire_6_15;
  wire [7:0] wire_6_16;
  wire [7:0] wire_6_17;
  wire [7:0] wire_6_18;
  assign wire_6 = wire_6_0|wire_6_1|wire_6_2|wire_6_3|wire_6_4|wire_6_5|wire_6_6|wire_6_7|wire_6_8|wire_6_9|wire_6_10|wire_6_11|wire_6_12|wire_6_13|wire_6_14|wire_6_15|wire_6_16|wire_6_17|wire_6_18;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [0:0] wire_10;
  wire [63:0] wire_11;
  wire [63:0] wire_11_0;
  wire [63:0] wire_11_1;
  wire [63:0] wire_11_2;
  wire [63:0] wire_11_3;
  wire [63:0] wire_11_4;
  wire [63:0] wire_11_5;
  wire [63:0] wire_11_6;
  wire [63:0] wire_11_7;
  wire [63:0] wire_11_8;
  wire [63:0] wire_11_9;
  wire [63:0] wire_11_10;
  wire [63:0] wire_11_11;
  wire [63:0] wire_11_12;
  wire [63:0] wire_11_13;
  wire [63:0] wire_11_14;
  wire [63:0] wire_11_15;
  wire [63:0] wire_11_16;
  wire [63:0] wire_11_17;
  assign wire_11 = wire_11_0|wire_11_1|wire_11_2|wire_11_3|wire_11_4|wire_11_5|wire_11_6|wire_11_7|wire_11_8|wire_11_9|wire_11_10|wire_11_11|wire_11_12|wire_11_13|wire_11_14|wire_11_15|wire_11_16|wire_11_17;
  wire [0:0] wire_12;
  wire [7:0] wire_13;
  wire [0:0] wire_14;
  wire [0:0] wire_15;
  wire [7:0] wire_16;
  wire [0:0] wire_17;
  wire [0:0] wire_18;
  wire [0:0] wire_19;
  wire [7:0] wire_20;
  wire [0:0] wire_21;
  wire [7:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [7:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [0:0] wire_31;
  wire [7:0] wire_32;
  wire [7:0] wire_32_0;
  wire [7:0] wire_32_1;
  wire [7:0] wire_32_2;
  wire [7:0] wire_32_3;
  wire [7:0] wire_32_4;
  wire [7:0] wire_32_5;
  wire [7:0] wire_32_6;
  wire [7:0] wire_32_7;
  wire [7:0] wire_32_8;
  wire [7:0] wire_32_9;
  wire [7:0] wire_32_10;
  wire [7:0] wire_32_11;
  wire [7:0] wire_32_12;
  wire [7:0] wire_32_13;
  wire [7:0] wire_32_14;
  assign wire_32 = wire_32_0|wire_32_1|wire_32_2|wire_32_3|wire_32_4|wire_32_5|wire_32_6|wire_32_7|wire_32_8|wire_32_9|wire_32_10|wire_32_11|wire_32_12|wire_32_13|wire_32_14;
  wire [0:0] wire_33;
  wire [0:0] wire_34;
  wire [0:0] wire_35;
  wire [0:0] wire_36;
  wire [0:0] wire_37;
  wire [7:0] wire_38;
  wire [7:0] wire_39;
  wire [7:0] wire_40;
  wire [7:0] wire_41;
  wire [0:0] wire_42;
  wire [0:0] wire_43;
  wire [7:0] wire_44;
  wire [0:0] wire_45;
  wire [0:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [7:0] wire_49;
  wire [0:0] wire_50;
  wire [0:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [63:0] wire_54;
  wire [15:0] wire_55;
  wire [7:0] wire_56;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [31:0] wire_62;
  wire [0:0] wire_63;
  wire [7:0] wire_64;
  wire [0:0] wire_65;
  wire [0:0] wire_66;
  wire [7:0] wire_67;
  wire [0:0] wire_68;
  wire [7:0] wire_69;
  wire [0:0] wire_70;
  wire [7:0] wire_71;
  wire [7:0] wire_72;
  wire [7:0] wire_73;
  wire [7:0] wire_74;
  wire [7:0] wire_75;
  wire [0:0] wire_76;
  wire [0:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [0:0] wire_80;
  wire [7:0] wire_81;
  wire [0:0] wire_82;
  wire [0:0] wire_83;
  wire [7:0] wire_84;
  wire [7:0] wire_85;
  wire [7:0] wire_85_0;
  wire [7:0] wire_85_1;
  assign wire_85 = wire_85_0|wire_85_1;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [0:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [7:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [7:0] wire_95;
  wire [0:0] wire_96;
  wire [0:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [7:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [0:0] wire_106;
  wire [0:0] wire_107;
  assign arch_output_enable = wire_107;
  wire [0:0] wire_108;
  wire [7:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [7:0] wire_114;
  wire [7:0] wire_115;
  wire [0:0] wire_116;
  wire [7:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [7:0] wire_121;
  wire [0:0] wire_122;
  wire [7:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;
  wire [7:0] wire_127;
  wire [0:0] wire_128;
  wire [0:0] wire_129;
  wire [0:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;
  wire [7:0] wire_133;
  wire [7:0] wire_133_0;
  wire [7:0] wire_133_1;
  wire [7:0] wire_133_2;
  assign wire_133 = wire_133_0|wire_133_1|wire_133_2;
  wire [0:0] wire_134;
  wire [0:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;
  wire [0:0] wire_138;
  wire [0:0] wire_139;
  wire [0:0] wire_140;
  wire [0:0] wire_140_0;
  wire [0:0] wire_140_1;
  wire [0:0] wire_140_2;
  wire [0:0] wire_140_3;
  wire [0:0] wire_140_4;
  wire [0:0] wire_140_5;
  wire [0:0] wire_140_6;
  wire [0:0] wire_140_7;
  assign wire_140 = wire_140_0|wire_140_1|wire_140_2|wire_140_3|wire_140_4|wire_140_5|wire_140_6|wire_140_7;
  wire [0:0] wire_141;
  wire [0:0] wire_142;
  wire [7:0] wire_143;
  wire [0:0] wire_144;
  wire [7:0] wire_145;
  wire [0:0] wire_146;
  wire [0:0] wire_147;
  wire [7:0] wire_148;
  wire [0:0] wire_149;
  wire [0:0] wire_150;
  wire [0:0] wire_151;
  wire [0:0] wire_152;
  wire [0:0] wire_153;
  wire [7:0] wire_154;
  wire [0:0] wire_155;
  wire [0:0] wire_156;
  wire [0:0] wire_157;
  wire [7:0] wire_158;
  wire [0:0] wire_159;
  wire [0:0] wire_160;
  wire [0:0] wire_161;
  wire [0:0] wire_162;
  wire [7:0] wire_163;
  wire [7:0] wire_164;
  wire [63:0] wire_165;
  wire [0:0] wire_166;
  wire [0:0] wire_167;
  wire [0:0] wire_168;
  wire [0:0] wire_169;
  wire [0:0] wire_170;
  wire [7:0] wire_171;
  wire [0:0] wire_172;
  wire [0:0] wire_173;
  wire [0:0] wire_174;
  wire [7:0] wire_175;
  wire [0:0] wire_176;
  wire [7:0] wire_177;
  wire [0:0] wire_178;
  wire [0:0] wire_179;
  wire [7:0] wire_180;
  wire [0:0] wire_181;
  wire [0:0] wire_182;
  wire [7:0] wire_183;
  wire [7:0] wire_184;
  wire [7:0] wire_184_0;
  wire [7:0] wire_184_1;
  assign wire_184 = wire_184_0|wire_184_1;
  wire [0:0] wire_185;
  wire [0:0] wire_186;
  wire [7:0] wire_187;
  wire [0:0] wire_188;
  wire [7:0] wire_189;
  wire [0:0] wire_190;
  wire [7:0] wire_191;
  wire [0:0] wire_192;
  wire [0:0] wire_193;
  wire [7:0] wire_194;
  wire [0:0] wire_195;
  wire [0:0] wire_196;
  wire [0:0] wire_197;
  wire [7:0] wire_198;
  wire [7:0] wire_198_0;
  wire [7:0] wire_198_1;
  assign wire_198 = wire_198_0|wire_198_1;
  wire [0:0] wire_199;
  wire [7:0] wire_200;
  wire [7:0] wire_201;
  wire [0:0] wire_202;
  wire [31:0] wire_203;
  wire [7:0] wire_204;
  wire [0:0] wire_205;
  wire [0:0] wire_206;
  wire [7:0] wire_207;
  wire [0:0] wire_208;
  wire [0:0] wire_209;
  wire [0:0] wire_210;
  wire [0:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [7:0] wire_214;
  wire [7:0] wire_214_0;
  wire [7:0] wire_214_1;
  assign wire_214 = wire_214_0|wire_214_1;
  wire [0:0] wire_215;
  wire [7:0] wire_216;
  wire [7:0] wire_217;
  wire [7:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [7:0] wire_221;
  wire [7:0] wire_221_0;
  wire [7:0] wire_221_1;
  assign wire_221 = wire_221_0|wire_221_1;
  wire [7:0] wire_222;
  wire [0:0] wire_223;
  wire [15:0] wire_224;
  wire [0:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [0:0] wire_228;
  wire [7:0] wire_229;
  wire [0:0] wire_230;
  wire [0:0] wire_231;
  wire [0:0] wire_232;
  wire [0:0] wire_233;
  wire [0:0] wire_234;
  wire [0:0] wire_235;
  wire [0:0] wire_236;
  wire [0:0] wire_237;
  wire [15:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [0:0] wire_242;
  wire [0:0] wire_243;
  wire [7:0] wire_244;
  wire [0:0] wire_245;
  wire [7:0] wire_246;
  wire [0:0] wire_247;
  wire [7:0] wire_248;
  wire [0:0] wire_249;
  wire [7:0] wire_250;
  wire [0:0] wire_251;
  wire [7:0] wire_252;
  wire [0:0] wire_253;
  wire [0:0] wire_254;
  wire [0:0] wire_255;
  wire [0:0] wire_256;
  wire [0:0] wire_257;
  wire [0:0] wire_258;
  wire [0:0] wire_259;
  wire [7:0] wire_260;
  wire [63:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [7:0] wire_265;
  wire [0:0] wire_266;
  wire [0:0] wire_267;
  wire [0:0] wire_268;
  wire [7:0] wire_269;
  wire [0:0] wire_270;
  wire [7:0] wire_271;
  wire [0:0] wire_272;
  wire [7:0] wire_273;
  wire [7:0] wire_274;
  wire [0:0] wire_275;
  wire [7:0] wire_276;
  wire [7:0] wire_277;
  wire [15:0] wire_278;
  wire [7:0] wire_279;
  wire [7:0] wire_280;
  wire [63:0] wire_281;
  wire [0:0] wire_282;
  wire [0:0] wire_283;
  wire [0:0] wire_284;
  wire [7:0] wire_285;
  wire [0:0] wire_286;
  wire [0:0] wire_287;
  wire [0:0] wire_288;
  wire [0:0] wire_289;
  wire [7:0] wire_290;
  wire [0:0] wire_291;
  wire [0:0] wire_292;
  wire [0:0] wire_293;
  wire [0:0] wire_294;
  wire [0:0] wire_295;
  wire [7:0] wire_296;
  wire [63:0] wire_297;
  wire [0:0] wire_298;
  wire [7:0] wire_299;
  wire [7:0] wire_300;
  wire [7:0] wire_301;
  wire [7:0] wire_302;
  wire [0:0] wire_303;
  wire [0:0] wire_304;
  wire [0:0] wire_305;
  wire [7:0] wire_306;
  wire [7:0] wire_307;
  wire [0:0] wire_308;

endmodule
