module Pixiez_Snake (clk, rst);
  parameter UUID = 0;
  parameter NAME = "";
  input wire clk;
  input wire rst;


  TC_Not # (.UUID(64'd680444558656414018 ^ UUID), .BIT_WIDTH(64'd1)) Not_0 (.in(wire_242), .out(wire_413));
  TC_Or3 # (.UUID(64'd534734424402985405 ^ UUID), .BIT_WIDTH(64'd1)) Or3_1 (.in0(wire_98), .in1(wire_442), .in2(wire_186), .out(wire_87));
  TC_Or3 # (.UUID(64'd4567130074526553310 ^ UUID), .BIT_WIDTH(64'd1)) Or3_2 (.in0(wire_52), .in1(wire_347), .in2(wire_228), .out(wire_250));
  TC_Or3 # (.UUID(64'd2737475285567390637 ^ UUID), .BIT_WIDTH(64'd1)) Or3_3 (.in0(wire_257), .in1(wire_133), .in2(wire_184), .out(wire_188));
  TC_Or3 # (.UUID(64'd1460121507051805330 ^ UUID), .BIT_WIDTH(64'd1)) Or3_4 (.in0(wire_188), .in1(wire_250), .in2(wire_67), .out(wire_229));
  TC_Not # (.UUID(64'd3263495404627770251 ^ UUID), .BIT_WIDTH(64'd1)) Not_5 (.in(wire_213), .out(wire_20));
  TC_DelayLine # (.UUID(64'd1861931133330004945 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_6 (.clk(clk), .rst(rst), .in(wire_20), .out(wire_213));
  TC_Not # (.UUID(64'd774824456586639901 ^ UUID), .BIT_WIDTH(64'd1)) Not_7 (.in(wire_263), .out(wire_455));
  TC_Or3 # (.UUID(64'd957665538453266802 ^ UUID), .BIT_WIDTH(64'd1)) Or3_8 (.in0(wire_146), .in1(wire_87), .in2(wire_143), .out(wire_263));
  TC_Add # (.UUID(64'd3301328818535174719 ^ UUID), .BIT_WIDTH(64'd8)) Add8_9 (.in0(wire_139), .in1(wire_80), .ci(wire_455), .out(wire_238), .co());
  TC_Or # (.UUID(64'd3186172645923730952 ^ UUID), .BIT_WIDTH(64'd1)) Or_10 (.in0(wire_372), .in1(wire_307), .out(wire_98));
  TC_Not # (.UUID(64'd4418713765798495162 ^ UUID), .BIT_WIDTH(64'd1)) Not_11 (.in(wire_4), .out(wire_318));
  TC_Or3 # (.UUID(64'd3359031826937924206 ^ UUID), .BIT_WIDTH(64'd1)) Or3_12 (.in0(wire_310), .in1(wire_338), .in2(wire_138), .out(wire_372));
  TC_Decoder3 # (.UUID(64'd4465221940936740645 ^ UUID)) Decoder3_13 (.dis(wire_60), .sel0(wire_158[0:0]), .sel1(wire_66[0:0]), .sel2(wire_261[0:0]), .out0(wire_52), .out1(wire_219), .out2(wire_187), .out3(wire_267), .out4(wire_89), .out5(wire_193), .out6(wire_138), .out7(wire_211));
  TC_Decoder3 # (.UUID(64'd664854618839101163 ^ UUID)) Decoder3_14 (.dis(wire_262), .sel0(wire_158[0:0]), .sel1(wire_66[0:0]), .sel2(wire_261[0:0]), .out0(wire_176), .out1(wire_228), .out2(wire_347), .out3(wire_291), .out4(wire_102), .out5(wire_204), .out6(wire_75), .out7(wire_331));
  TC_Decoder3 # (.UUID(64'd388458847481545701 ^ UUID)) Decoder3_15 (.dis(wire_407), .sel0(wire_158[0:0]), .sel1(wire_66[0:0]), .sel2(wire_261[0:0]), .out0(wire_285), .out1(wire_28), .out2(wire_345), .out3(wire_220), .out4(wire_166), .out5(wire_6), .out6(wire_179), .out7(wire_104));
  TC_Decoder3 # (.UUID(64'd1325274093033025990 ^ UUID)) Decoder3_16 (.dis(wire_48), .sel0(wire_158[0:0]), .sel1(wire_66[0:0]), .sel2(wire_261[0:0]), .out0(wire_402), .out1(wire_184), .out2(wire_133), .out3(wire_257), .out4(wire_68), .out5(wire_118), .out6(wire_25), .out7(wire_371));
  TC_Not # (.UUID(64'd56215910927289989 ^ UUID), .BIT_WIDTH(64'd1)) Not_17 (.in(wire_412), .out(wire_60));
  TC_Not # (.UUID(64'd1568445558185814797 ^ UUID), .BIT_WIDTH(64'd1)) Not_18 (.in(wire_449), .out(wire_48));
  TC_Not # (.UUID(64'd3688819333690076749 ^ UUID), .BIT_WIDTH(64'd1)) Not_19 (.in(wire_180), .out(wire_407));
  TC_Not # (.UUID(64'd2914649659429896514 ^ UUID), .BIT_WIDTH(64'd1)) Not_20 (.in(wire_474), .out(wire_262));
  TC_Maker8 # (.UUID(64'd4274226248529413390 ^ UUID)) Maker8_21 (.in0(wire_52), .in1(wire_219), .in2(wire_187), .in3(wire_267), .in4(wire_89), .in5(wire_193), .in6(wire_138), .in7(wire_211), .out(wire_201));
  TC_Maker8 # (.UUID(64'd2503620967526902392 ^ UUID)) Maker8_22 (.in0(wire_176), .in1(wire_228), .in2(wire_347), .in3(wire_291), .in4(wire_102), .in5(wire_204), .in6(wire_75), .in7(wire_331), .out(wire_129));
  TC_Maker8 # (.UUID(64'd736697256551715288 ^ UUID)) Maker8_23 (.in0(wire_285), .in1(wire_28), .in2(wire_345), .in3(wire_220), .in4(wire_166), .in5(wire_6), .in6(wire_179), .in7(wire_104), .out(wire_175));
  TC_Maker8 # (.UUID(64'd832968618284013991 ^ UUID)) Maker8_24 (.in0(wire_402), .in1(wire_184), .in2(wire_133), .in3(wire_257), .in4(wire_68), .in5(wire_118), .in6(wire_25), .in7(wire_371), .out(wire_202));
  TC_Or3 # (.UUID(64'd2334335797361251671 ^ UUID), .BIT_WIDTH(64'd1)) Or3_25 (.in0(wire_75), .in1(wire_331), .in2(wire_267), .out(wire_338));
  TC_Or3 # (.UUID(64'd4505646521355499044 ^ UUID), .BIT_WIDTH(64'd1)) Or3_26 (.in0(wire_118), .in1(wire_371), .in2(wire_285), .out(wire_307));
  TC_Or3 # (.UUID(64'd2771484508194729184 ^ UUID), .BIT_WIDTH(64'd1)) Or3_27 (.in0(wire_6), .in1(wire_166), .in2(wire_220), .out(wire_41));
  TC_Or3 # (.UUID(64'd2848731522163985212 ^ UUID), .BIT_WIDTH(64'd1)) Or3_28 (.in0(wire_176), .in1(wire_104), .in2(wire_179), .out(wire_383));
  TC_DelayLine # (.UUID(64'd1068115119822942229 ^ UUID), .BIT_WIDTH(64'd8)) DelayLine8_29 (.clk(clk), .rst(rst), .in(wire_13[7:0]), .out(wire_424));
  TC_DelayLine # (.UUID(64'd804044612046236745 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_30 (.clk(clk), .rst(rst), .in(wire_336), .out(wire_242));
  TC_Splitter16 # (.UUID(64'd1875228578544666958 ^ UUID)) Splitter16_31 (.in(wire_357), .out0(wire_456), .out1(wire_260));
  TC_Maker16 # (.UUID(64'd3608744494562313405 ^ UUID)) Maker16_32 (.in0({{7{1'b0}}, wire_413 }), .in1(wire_436), .out(wire_357));
  TC_Or3 # (.UUID(64'd3746619389515595809 ^ UUID), .BIT_WIDTH(64'd1)) Or3_33 (.in0(wire_29), .in1(wire_72), .in2(wire_366), .out(wire_336));
  TC_Not # (.UUID(64'd966737772035534885 ^ UUID), .BIT_WIDTH(64'd1)) Not_34 (.in(wire_254[0:0]), .out(wire_444));
  TC_Not # (.UUID(64'd424140961992658426 ^ UUID), .BIT_WIDTH(64'd1)) Not_35 (.in(wire_10[0:0]), .out(wire_459));
  TC_Splitter32 # (.UUID(64'd2809680451032690949 ^ UUID)) Splitter32_36 (.in(wire_69), .out0(wire_358), .out1(), .out2(), .out3());
  TC_Constant # (.UUID(64'd2117984546099265654 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_37 (.out(wire_295));
  TC_Mux # (.UUID(64'd2353982102422779838 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_38 (.sel(wire_274), .in0(wire_0), .in1(wire_295), .out(wire_411));
  TC_Add # (.UUID(64'd4134817076244850895 ^ UUID), .BIT_WIDTH(64'd8)) Add8_39 (.in0(wire_2), .in1(wire_411), .ci(1'd0), .out(wire_340), .co());
  TC_Constant # (.UUID(64'd1952156418708934468 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_40 (.out(wire_258));
  TC_Mux # (.UUID(64'd4094225513381061300 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_41 (.sel(wire_205), .in0(wire_0), .in1(wire_258), .out(wire_364));
  TC_Neg # (.UUID(64'd102576365000716770 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_42 (.in(wire_364), .out(wire_135));
  TC_Add # (.UUID(64'd2689942381287690498 ^ UUID), .BIT_WIDTH(64'd8)) Add8_43 (.in0(wire_2), .in1(wire_135), .ci(1'd0), .out(wire_252), .co());
  TC_Mul # (.UUID(64'd3289678684259179587 ^ UUID), .BIT_WIDTH(64'd8)) Mul8_44 (.in0(wire_2), .in1(wire_0), .out0(wire_57), .out1());
  TC_Switch # (.UUID(64'd3227644779488857845 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_45 (.en(wire_154), .in(wire_57), .out(wire_13_11[7:0]));
  TC_Switch # (.UUID(64'd4137287338459891824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_46 (.en(wire_40), .in(wire_252), .out(wire_13_13[7:0]));
  TC_Switch # (.UUID(64'd1351346083360514605 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_47 (.en(wire_105), .in(wire_340), .out(wire_13_15[7:0]));
  TC_Splitter8 # (.UUID(64'd4357406098891943912 ^ UUID)) Splitter8_48 (.in(wire_358), .out0(wire_296), .out1(wire_100), .out2(wire_154), .out3(wire_79), .out4(wire_170), .out5(wire_274), .out6(wire_205), .out7(wire_293));
  TC_Not # (.UUID(64'd3532098913873322011 ^ UUID), .BIT_WIDTH(64'd1)) Not_49 (.in(wire_287[0:0]), .out(wire_290));
  TC_Switch # (.UUID(64'd2937048381182156076 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_50 (.en(wire_4), .in(wire_230), .out(wire_2_2));
  TC_Switch # (.UUID(64'd412107824868226985 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_51 (.en(wire_318), .in(wire_230), .out(wire_127));
  TC_Switch # (.UUID(64'd1458121506772114657 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_52 (.en(wire_254[0:0]), .in(wire_270), .out(wire_0_2));
  TC_Switch # (.UUID(64'd2507210810598866832 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_53 (.en(wire_444), .in(wire_270), .out(wire_130));
  TC_Switch # (.UUID(64'd1855204595012977435 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_54 (.en(wire_287[0:0]), .in(wire_63), .out(wire_13_8[7:0]));
  TC_Switch # (.UUID(64'd1879885438156656135 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_55 (.en(wire_290), .in(wire_63), .out(wire_203));
  TC_Splitter16 # (.UUID(64'd4592662178931061204 ^ UUID)) Splitter16_56 (.in(wire_214), .out0(wire_88), .out1(wire_10));
  TC_Or3 # (.UUID(64'd1577578265915915529 ^ UUID), .BIT_WIDTH(64'd1)) Or3_57 (.in0(wire_88[0:0]), .in1(wire_10[0:0]), .in2(wire_146), .out(wire_73));
  TC_Switch # (.UUID(64'd2610614871112416436 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_58 (.en(wire_88[0:0]), .in(wire_414[7:0]), .out(wire_160));
  TC_Switch # (.UUID(64'd165300680693317419 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_59 (.en(wire_88[0:0]), .in(wire_91[7:0]), .out(wire_270));
  TC_Switch # (.UUID(64'd2260740780324363689 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_60 (.en(wire_73), .in(wire_106[7:0]), .out(wire_230));
  TC_Mux # (.UUID(64'd4528590367296190010 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_61 (.sel(wire_459), .in0(wire_91[7:0]), .in1(wire_160), .out(wire_63));
  TC_Splitter16 # (.UUID(64'd2701914707745210702 ^ UUID)) Splitter16_62 (.in(wire_344), .out0(wire_287), .out1(wire_254));
  TC_Maker16 # (.UUID(64'd1365218859602849489 ^ UUID)) Maker16_63 (.in0({{7{1'b0}}, wire_370 }), .in1({{7{1'b0}}, wire_420 }), .out(wire_344));
  TC_Switch # (.UUID(64'd2155635750972134594 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_64 (.en(wire_242), .in(wire_424), .out(wire_436));
  TC_Mux # (.UUID(64'd1791751815309933921 ^ UUID), .BIT_WIDTH(64'd8)) Mux8_65 (.sel(wire_456[0:0]), .in0(wire_260), .in1(wire_34), .out(wire_139));
  TC_Maker16 # (.UUID(64'd3395313277560932739 ^ UUID)) Maker16_66 (.in0({{7{1'b0}}, wire_143 }), .in1({{7{1'b0}}, wire_87 }), .out(wire_214));
  TC_Not # (.UUID(64'd3453103485371531751 ^ UUID), .BIT_WIDTH(64'd1)) Not_67 (.in(wire_20), .out(wire_82));
  TC_Counter # (.UUID(64'd1171561396707692790 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_68 (.clk(clk), .rst(rst), .save(wire_20), .in(wire_238), .out(wire_415));
  TC_Counter # (.UUID(64'd2621291279726673638 ^ UUID), .BIT_WIDTH(64'd8), .count(8'd1)) Counter8_69 (.clk(clk), .rst(rst), .save(wire_213), .in(wire_238), .out(wire_392));
  TC_Switch # (.UUID(64'd1839974249620431880 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_70 (.en(wire_82), .in(wire_415), .out(wire_34_0));
  TC_Switch # (.UUID(64'd1170108399670313272 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_71 (.en(wire_20), .in(wire_392), .out(wire_34_1));
  TC_Constant # (.UUID(64'd358007510611002277 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h2)) Constant8_72 (.out(wire_428));
  TC_Constant # (.UUID(64'd3874548421935569254 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h3)) Constant8_73 (.out(wire_453));
  TC_Constant # (.UUID(64'd1203375723678859801 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h4)) Constant8_74 (.out(wire_389));
  TC_Switch # (.UUID(64'd1933124139798812111 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_75 (.en(wire_146), .in(wire_428), .out(wire_80_2));
  TC_Switch # (.UUID(64'd287643768980040071 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_76 (.en(wire_87), .in(wire_453), .out(wire_80_1));
  TC_Switch # (.UUID(64'd4195386940103341620 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_77 (.en(wire_143), .in(wire_389), .out(wire_80_0));
  TC_Splitter8 # (.UUID(64'd2599557092287595297 ^ UUID)) Splitter8_78 (.in(wire_5[7:0]), .out0(wire_112), .out1(wire_445), .out2(wire_452), .out3(wire_467), .out4(wire_401), .out5(wire_370), .out6(wire_420), .out7(wire_4));
  TC_Ram # (.UUID(64'd1708105537810654235 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd256)) Ram_79 (.clk(clk), .rst(rst), .load(wire_7), .save(wire_353), .address({{24{1'b0}}, wire_0 }), .in0({{56{1'b0}}, wire_2 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_13_0), .out1(), .out2(), .out3());
  TC_Ram # (.UUID(64'd97660009947370162 ^ UUID), .WORD_WIDTH(64'd16), .WORD_COUNT(64'd128)) Ram_80 (.clk(clk), .rst(rst), .load(wire_162), .save(wire_22), .address({{24{1'b0}}, wire_297 }), .in0({{56{1'b0}}, wire_238 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_181), .out1(), .out2(), .out3());
  TC_Or # (.UUID(64'd733084299857471502 ^ UUID), .BIT_WIDTH(64'd1)) Or_81 (.in0(wire_22), .in1(wire_162), .out(wire_29));
  TC_Splitter32 # (.UUID(64'd3048987527585864498 ^ UUID)) Splitter32_82 (.in(wire_69), .out0(), .out1(wire_167), .out2(), .out3(wire_327));
  TC_Or # (.UUID(64'd4064324485441264957 ^ UUID), .BIT_WIDTH(64'd1)) Or_83 (.in0(wire_162), .in1(wire_22), .out(wire_314));
  TC_Switch # (.UUID(64'd2955305895674404779 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_84 (.en(wire_162), .in(wire_181[7:0]), .out(wire_13_4[7:0]));
  TC_Switch # (.UUID(64'd3592902196704226444 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_85 (.en(wire_22), .in(wire_2), .out(wire_13_3[7:0]));
  TC_Register # (.UUID(64'd4471884361578131577 ^ UUID), .BIT_WIDTH(64'd8)) Register8_86 (.clk(clk), .rst(rst), .load(wire_314), .save(wire_314), .in(wire_168), .out(wire_12));
  TC_Switch # (.UUID(64'd4562232227874677430 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_87 (.en(wire_22), .in(wire_231), .out(wire_168_0));
  TC_Switch # (.UUID(64'd114510401986147547 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_88 (.en(wire_22), .in(wire_168), .out(wire_297_0));
  TC_Add # (.UUID(64'd263770477141513169 ^ UUID), .BIT_WIDTH(64'd8)) Add8_89 (.in0(wire_46), .in1(wire_12), .ci(1'd0), .out(wire_231), .co());
  TC_Switch # (.UUID(64'd2865125256828769888 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_90 (.en(wire_162), .in(wire_386), .out(wire_168_1));
  TC_Switch # (.UUID(64'd1945149825988830027 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_91 (.en(wire_162), .in(wire_12), .out(wire_297_1));
  TC_Constant # (.UUID(64'd2864754851009931669 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_92 (.out(wire_46));
  TC_Neg # (.UUID(64'd1766191137768834313 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_93 (.in(wire_46), .out(wire_475));
  TC_Add # (.UUID(64'd1197352873015043648 ^ UUID), .BIT_WIDTH(64'd8)) Add8_94 (.in0(wire_12), .in1(wire_475), .ci(1'd0), .out(wire_386), .co());
  TC_Splitter8 # (.UUID(64'd3473615707126412287 ^ UUID)) Splitter8_95 (.in(wire_327), .out0(wire_353), .out1(wire_7), .out2(), .out3(), .out4(), .out5(), .out6(), .out7(wire_126));
  TC_Constant # (.UUID(64'd3007591360524826255 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h0)) Constant8_96 (.out(wire_273));
  TC_Or # (.UUID(64'd3353986015329929110 ^ UUID), .BIT_WIDTH(64'd1)) Or_97 (.in0(wire_56), .in1(wire_172), .out(wire_217));
  TC_LessU # (.UUID(64'd2857803572762207218 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_98 (.in0(wire_0), .in1(wire_2), .out(wire_172));
  TC_Not # (.UUID(64'd3713135576456282771 ^ UUID), .BIT_WIDTH(64'd1)) Not_99 (.in(wire_56), .out(wire_223));
  TC_Or # (.UUID(64'd1283831029887634373 ^ UUID), .BIT_WIDTH(64'd1)) Or_100 (.in0(wire_14), .in1(wire_56), .out(wire_320));
  TC_Equal # (.UUID(64'd3249866343864622854 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_101 (.in0(wire_2), .in1(wire_0), .out(wire_56));
  TC_LessU # (.UUID(64'd2949327424893302673 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_102 (.in0(wire_2), .in1(wire_0), .out(wire_14));
  TC_Equal # (.UUID(64'd3467215832225421993 ^ UUID), .BIT_WIDTH(64'd8)) Equal8_103 (.in0(wire_273), .in1(wire_2), .out(wire_451));
  TC_Constant # (.UUID(64'd4251321236624205294 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_104 (.out(wire_440));
  TC_Switch # (.UUID(64'd4268044874154730043 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_105 (.en(wire_194), .in(wire_440), .out(wire_72_7));
  TC_Switch # (.UUID(64'd1386783397630713083 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_106 (.en(wire_207), .in(wire_451), .out(wire_72_5));
  TC_Switch # (.UUID(64'd1155028069485320511 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_107 (.en(wire_315), .in(wire_14), .out(wire_72_3));
  TC_Switch # (.UUID(64'd3348470806054818924 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_108 (.en(wire_245), .in(wire_320), .out(wire_72_0));
  TC_Switch # (.UUID(64'd1041869814803847902 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_109 (.en(wire_147), .in(wire_56), .out(wire_72_1));
  TC_Switch # (.UUID(64'd4055918702281020749 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_110 (.en(wire_178), .in(wire_223), .out(wire_72_2));
  TC_Switch # (.UUID(64'd3083535767069260986 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_111 (.en(wire_39), .in(wire_217), .out(wire_72_4));
  TC_Switch # (.UUID(64'd2913504031160566908 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_112 (.en(wire_49), .in(wire_172), .out(wire_72_6));
  TC_Splitter8 # (.UUID(64'd1194059391229914692 ^ UUID)) Splitter8_113 (.in(wire_167), .out0(wire_194), .out1(wire_207), .out2(wire_315), .out3(wire_245), .out4(wire_147), .out5(wire_178), .out6(wire_39), .out7(wire_49));
  TC_Register # (.UUID(64'd1786549938381629068 ^ UUID), .BIT_WIDTH(64'd8)) Register8_114 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_375), .in(wire_13[7:0]), .out(wire_319));
  TC_Register # (.UUID(64'd2601905860340903537 ^ UUID), .BIT_WIDTH(64'd8)) Register8_115 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_341), .in(wire_13[7:0]), .out(wire_346));
  TC_Register # (.UUID(64'd2818150811460271121 ^ UUID), .BIT_WIDTH(64'd8)) Register8_116 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_351), .in(wire_13[7:0]), .out(wire_37));
  TC_Register # (.UUID(64'd3810474016475870525 ^ UUID), .BIT_WIDTH(64'd8)) Register8_117 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_173), .in(wire_13[7:0]), .out(wire_15));
  TC_Register # (.UUID(64'd1636002980180907684 ^ UUID), .BIT_WIDTH(64'd8)) Register8_118 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_417), .in(wire_13[7:0]), .out(wire_356));
  TC_Register # (.UUID(64'd3256658416273011892 ^ UUID), .BIT_WIDTH(64'd8)) Register8_119 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_391), .in(wire_13[7:0]), .out(wire_152));
  TC_Register # (.UUID(64'd2526494128293687363 ^ UUID), .BIT_WIDTH(64'd8)) Register8_120 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_443), .in(wire_13[7:0]), .out(wire_190));
  TC_Register # (.UUID(64'd3472073544120575095 ^ UUID), .BIT_WIDTH(64'd8)) Register8_121 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_150), .in(wire_13[7:0]), .out(wire_311));
  TC_Register # (.UUID(64'd542285582491664182 ^ UUID), .BIT_WIDTH(64'd8)) Register8_122 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_233), .in(wire_13[7:0]), .out(wire_43));
  TC_Register # (.UUID(64'd2124618488310653916 ^ UUID), .BIT_WIDTH(64'd8)) Register8_123 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_374), .in(wire_13[7:0]), .out(wire_208));
  TC_Register # (.UUID(64'd240222191994770064 ^ UUID), .BIT_WIDTH(64'd8)) Register8_124 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_90), .in(wire_13[7:0]), .out(wire_313));
  TC_Switch # (.UUID(64'd2919893529833212573 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_125 (.en(wire_337), .in(wire_37), .out(wire_2_18));
  TC_Switch # (.UUID(64'd2892052628952263194 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_126 (.en(wire_410), .in(wire_37), .out(wire_0_18));
  TC_Switch # (.UUID(64'd1045466942081498185 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_127 (.en(wire_218), .in(wire_15), .out(wire_2_17));
  TC_Switch # (.UUID(64'd4352568465751771503 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_128 (.en(wire_93), .in(wire_15), .out(wire_0_17));
  TC_Switch # (.UUID(64'd294837876173931186 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_129 (.en(wire_335), .in(wire_190), .out(wire_2_16));
  TC_Switch # (.UUID(64'd718804107324007425 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_130 (.en(wire_276), .in(wire_190), .out(wire_0_16));
  TC_Switch # (.UUID(64'd2106337721725300490 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_131 (.en(wire_169), .in(wire_43), .out(wire_2_15));
  TC_Switch # (.UUID(64'd1382626067278158580 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_132 (.en(wire_199), .in(wire_43), .out(wire_0_15));
  TC_Switch # (.UUID(64'd4280389427710179554 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_133 (.en(wire_119), .in(wire_311), .out(wire_2_14));
  TC_Switch # (.UUID(64'd2870197787210989981 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_134 (.en(wire_246), .in(wire_311), .out(wire_0_14));
  TC_Switch # (.UUID(64'd1025076596807518358 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_135 (.en(wire_423), .in(wire_356), .out(wire_2_13));
  TC_Switch # (.UUID(64'd961920732700576390 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_136 (.en(wire_419), .in(wire_356), .out(wire_0_13));
  TC_Switch # (.UUID(64'd455633754159767112 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_137 (.en(wire_18), .in(wire_208), .out(wire_2_12));
  TC_Switch # (.UUID(64'd3572372897415253218 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_138 (.en(wire_447), .in(wire_208), .out(wire_0_12));
  TC_Switch # (.UUID(64'd2693638907193452534 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_139 (.en(wire_235), .in(wire_152), .out(wire_2_11));
  TC_Switch # (.UUID(64'd4344217990313000347 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_140 (.en(wire_395), .in(wire_152), .out(wire_0_11));
  TC_Switch # (.UUID(64'd258289412669476303 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_141 (.en(wire_103), .in(wire_346), .out(wire_2_10));
  TC_Switch # (.UUID(64'd4506884556720173301 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_142 (.en(wire_405), .in(wire_346), .out(wire_0_10));
  TC_Switch # (.UUID(64'd3160999002775359256 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_143 (.en(wire_281), .in(wire_319), .out(wire_2_9));
  TC_Switch # (.UUID(64'd4258632307214665985 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_144 (.en(wire_253), .in(wire_319), .out(wire_0_9));
  TC_Switch # (.UUID(64'd1115547685276398812 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_145 (.en(wire_171), .in(wire_313), .out(wire_2_8));
  TC_Switch # (.UUID(64'd2594916914153554215 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_146 (.en(wire_454), .in(wire_313), .out(wire_0_8));
  TC_Switch # (.UUID(64'd2067768058777429209 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_147 (.en(wire_342), .in(wire_323), .out(wire_0_6));
  TC_Switch # (.UUID(64'd1049797112137663963 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_148 (.en(wire_123), .in(wire_323), .out(wire_2_4));
  TC_Switch # (.UUID(64'd4067917907888700042 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_149 (.en(wire_249), .in(wire_280), .out(wire_0_7));
  TC_Switch # (.UUID(64'd3311537942366866912 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_150 (.en(wire_422), .in(wire_280), .out(wire_2_7));
  TC_Register # (.UUID(64'd1377807017811864986 ^ UUID), .BIT_WIDTH(64'd8)) Register8_151 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_221), .in(wire_13[7:0]), .out(wire_280));
  TC_Register # (.UUID(64'd1236368519178447850 ^ UUID), .BIT_WIDTH(64'd8)) Register8_152 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_301), .in(wire_13[7:0]), .out(wire_323));
  TC_Splitter8 # (.UUID(64'd2271575679199078636 ^ UUID)) Splitter8_153 (.in(wire_328), .out0(), .out1(), .out2(wire_92), .out3(wire_151), .out4(wire_22), .out5(wire_162), .out6(), .out7());
  TC_Splitter32 # (.UUID(64'd261396410293330702 ^ UUID)) Splitter32_154 (.in(wire_69), .out0(), .out1(), .out2(), .out3(wire_328));
  TC_Ram # (.UUID(64'd4117401978527469154 ^ UUID), .WORD_WIDTH(64'd8), .WORD_COUNT(64'd32)) Ram_155 (.clk(clk), .rst(rst), .load(wire_151), .save(wire_92), .address({{24{1'b0}}, wire_128 }), .in0({{56{1'b0}}, wire_2 }), .in1(64'd0), .in2(64'd0), .in3(64'd0), .out0(wire_13_2), .out1(), .out2(), .out3());
  TC_Switch # (.UUID(64'd3226929204346999104 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_156 (.en(wire_79), .in({{7{1'b0}}, wire_393 }), .out(wire_13_7[7:0]));
  TC_Switch # (.UUID(64'd3161290829479641019 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_157 (.en(wire_170), .in(wire_446), .out(wire_13_6[7:0]));
  TC_Switch # (.UUID(64'd3115314308242652354 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_158 (.en(wire_293), .in(wire_406), .out(wire_13_5[7:0]));
  TC_Neg # (.UUID(64'd77226668367061539 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_159 (.in(wire_2), .out(wire_446));
  TC_Or # (.UUID(64'd1380170131908116772 ^ UUID), .BIT_WIDTH(64'd1)) Or_160 (.in0(wire_205), .in1(wire_100), .out(wire_40));
  TC_Constant # (.UUID(64'd4166492318356521758 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_161 (.out(wire_17));
  TC_Constant # (.UUID(64'd1678158762324492118 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_162 (.out(wire_237));
  TC_Ashr # (.UUID(64'd1558764338386234982 ^ UUID), .BIT_WIDTH(64'd8)) Ashr8_163 (.in(wire_2), .shift(wire_237), .out(wire_406));
  TC_Constant # (.UUID(64'd2997253212554120558 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_164 (.out(wire_3));
  TC_Constant # (.UUID(64'd3797620182831446698 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h1)) Constant8_165 (.out(wire_283));
  TC_Neg # (.UUID(64'd3558537661740369771 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_166 (.in(wire_283), .out(wire_479));
  TC_Register # (.UUID(64'd2759537605007938592 ^ UUID), .BIT_WIDTH(64'd8)) Register8_167 (.clk(clk), .rst(rst), .load(wire_210), .save(wire_210), .in(wire_215), .out(wire_19));
  TC_Switch # (.UUID(64'd929829793202303828 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_168 (.en(wire_92), .in(wire_466), .out(wire_215_0));
  TC_Switch # (.UUID(64'd3728124673178845213 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_169 (.en(wire_92), .in(wire_215), .out(wire_128_1));
  TC_Add # (.UUID(64'd1902099203606853874 ^ UUID), .BIT_WIDTH(64'd8)) Add8_170 (.in0(wire_283), .in1(wire_19), .ci(1'd0), .out(wire_466), .co());
  TC_Switch # (.UUID(64'd3498208789273416986 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_171 (.en(wire_151), .in(wire_142), .out(wire_215_1));
  TC_Switch # (.UUID(64'd1321154288873073244 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_172 (.en(wire_151), .in(wire_19), .out(wire_128_0));
  TC_Or # (.UUID(64'd1321825518205599775 ^ UUID), .BIT_WIDTH(64'd1)) Or_173 (.in0(wire_151), .in1(wire_92), .out(wire_210));
  TC_Add # (.UUID(64'd4199771119303044950 ^ UUID), .BIT_WIDTH(64'd8)) Add8_174 (.in0(wire_19), .in1(wire_479), .ci(1'd0), .out(wire_142), .co());
  TC_Switch # (.UUID(64'd81193405753331740 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_175 (.en(wire_394), .in(wire_317), .out(wire_13_19[7:0]));
  TC_Switch # (.UUID(64'd4415608983622849585 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_176 (.en(wire_33), .in(wire_189), .out(wire_13_18[7:0]));
  TC_And # (.UUID(64'd1669263777784106749 ^ UUID), .BIT_WIDTH(64'd8)) And8_177 (.in0(wire_2), .in1(wire_0), .out(wire_317));
  TC_Or # (.UUID(64'd873622160744398625 ^ UUID), .BIT_WIDTH(64'd8)) Or8_178 (.in0(wire_2), .in1(wire_0), .out(wire_189));
  TC_Xor # (.UUID(64'd2690694932656199993 ^ UUID), .BIT_WIDTH(64'd8)) Xor8_179 (.in0(wire_2), .in1(wire_0), .out(wire_312));
  TC_Not # (.UUID(64'd3218967706620565239 ^ UUID), .BIT_WIDTH(64'd8)) Not8_180 (.in(wire_2), .out(wire_477));
  TC_Shl # (.UUID(64'd3160996752802486419 ^ UUID), .BIT_WIDTH(64'd8)) Shl8_181 (.in(wire_2), .shift(wire_17), .out(wire_399));
  TC_Shr # (.UUID(64'd1938059414175291844 ^ UUID), .BIT_WIDTH(64'd8)) Shr8_182 (.in(wire_2), .shift(wire_17), .out(wire_116));
  TC_Rol # (.UUID(64'd379560068498716864 ^ UUID), .BIT_WIDTH(64'd8)) Rol8_183 (.in(wire_2), .shift(wire_17), .out(wire_367));
  TC_Ror # (.UUID(64'd4299448326393726552 ^ UUID), .BIT_WIDTH(64'd8)) Ror8_184 (.in(wire_2), .shift(wire_17), .out(wire_282));
  TC_Switch # (.UUID(64'd2309803132069263134 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_185 (.en(wire_251), .in(wire_312), .out(wire_13_17[7:0]));
  TC_Switch # (.UUID(64'd2923996340214116429 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_186 (.en(wire_334), .in(wire_477), .out(wire_13_16[7:0]));
  TC_Switch # (.UUID(64'd2407013580594625997 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_187 (.en(wire_247), .in(wire_116), .out(wire_13_14[7:0]));
  TC_Switch # (.UUID(64'd3621734594009664278 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_188 (.en(wire_302), .in(wire_399), .out(wire_13_12[7:0]));
  TC_Switch # (.UUID(64'd1878036650580289106 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_189 (.en(wire_196), .in(wire_282), .out(wire_13_9[7:0]));
  TC_Switch # (.UUID(64'd4077902765271428258 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_190 (.en(wire_377), .in(wire_367), .out(wire_13_10[7:0]));
  TC_Splitter8 # (.UUID(64'd772965213957027290 ^ UUID)) Splitter8_191 (.in(wire_448), .out0(wire_394), .out1(wire_33), .out2(wire_251), .out3(wire_334), .out4(wire_247), .out5(wire_302), .out6(wire_196), .out7(wire_377));
  TC_Splitter32 # (.UUID(64'd3454244281776476436 ^ UUID)) Splitter32_192 (.in(wire_69), .out0(), .out1(), .out2(wire_448), .out3());
  TC_Register # (.UUID(64'd1044465739269958273 ^ UUID), .BIT_WIDTH(64'd8)) Register8_193 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_232), .in(wire_13[7:0]), .out(wire_97));
  TC_Register # (.UUID(64'd1014775350705063680 ^ UUID), .BIT_WIDTH(64'd8)) Register8_194 (.clk(clk), .rst(rst), .load(wire_3), .save(wire_206), .in(wire_13[7:0]), .out(wire_161));
  TC_Switch # (.UUID(64'd17400449972985902 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_195 (.en(wire_53), .in(wire_161), .out(wire_2_3));
  TC_Switch # (.UUID(64'd1757317349619379473 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_196 (.en(wire_373), .in(wire_161), .out(wire_0_3));
  TC_Switch # (.UUID(64'd347935731390232235 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_197 (.en(wire_306), .in(wire_97), .out(wire_2_1));
  TC_Switch # (.UUID(64'd347572746678109137 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_198 (.en(wire_387), .in(wire_97), .out(wire_0_1));
  TC_Switch # (.UUID(64'd117201099522242557 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_199 (.en(wire_185), .in(wire_238), .out(wire_2_0));
  TC_Switch # (.UUID(64'd1134152020965279556 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_200 (.en(wire_461), .in(wire_238), .out(wire_0_0));
  TC_Not # (.UUID(64'd2075639373923651350 ^ UUID), .BIT_WIDTH(64'd1)) Not_201 (.in(wire_113), .out(wire_390));
  TC_And # (.UUID(64'd754894496948066040 ^ UUID), .BIT_WIDTH(64'd1)) And_202 (.in0(wire_113), .in1(wire_125), .out(wire_144));
  TC_Or # (.UUID(64'd805549193662201184 ^ UUID), .BIT_WIDTH(64'd1)) Or_203 (.in0(wire_125), .in1(wire_390), .out(wire_85));
  TC_Decoder3 # (.UUID(64'd3761069498695685674 ^ UUID)) Decoder3_204 (.dis(wire_115), .sel0(wire_244), .sel1(wire_225), .sel2(wire_74), .out0(wire_337), .out1(wire_218), .out2(wire_335), .out3(wire_169), .out4(wire_119), .out5(wire_423), .out6(wire_18), .out7(wire_235));
  TC_Decoder3 # (.UUID(64'd1604216519862450208 ^ UUID)) Decoder3_205 (.dis(wire_85), .sel0(wire_244), .sel1(wire_225), .sel2(wire_74), .out0(wire_103), .out1(wire_281), .out2(wire_171), .out3(wire_422), .out4(wire_123), .out5(wire_53), .out6(wire_306), .out7(wire_27));
  TC_Or # (.UUID(64'd259192617280007518 ^ UUID), .BIT_WIDTH(64'd1)) Or_206 (.in0(wire_86), .in1(wire_480), .out(wire_71));
  TC_Decoder3 # (.UUID(64'd1295781503081853777 ^ UUID)) Decoder3_207 (.dis(wire_458), .sel0(wire_47), .sel1(wire_155), .sel2(wire_275), .out0(wire_410), .out1(wire_93), .out2(wire_276), .out3(wire_199), .out4(wire_246), .out5(wire_419), .out6(wire_447), .out7(wire_395));
  TC_Decoder3 # (.UUID(64'd57268074239693712 ^ UUID)) Decoder3_208 (.dis(wire_71), .sel0(wire_47), .sel1(wire_155), .sel2(wire_275), .out0(wire_405), .out1(wire_253), .out2(wire_454), .out3(wire_249), .out4(wire_342), .out5(wire_373), .out6(wire_387), .out7(wire_265));
  TC_Or # (.UUID(64'd1404831056388826959 ^ UUID), .BIT_WIDTH(64'd1)) Or_209 (.in0(wire_95), .in1(wire_145), .out(wire_94));
  TC_And # (.UUID(64'd2552562799264486541 ^ UUID), .BIT_WIDTH(64'd1)) And_210 (.in0(wire_240), .in1(wire_95), .out(wire_65));
  TC_Decoder3 # (.UUID(64'd762150619108810778 ^ UUID)) Decoder3_211 (.dis(wire_94), .sel0(wire_136), .sel1(wire_21), .sel2(wire_329), .out0(wire_341), .out1(wire_375), .out2(wire_90), .out3(wire_221), .out4(wire_301), .out5(wire_206), .out6(wire_232), .out7());
  TC_Decoder3 # (.UUID(64'd494457670381439667 ^ UUID)) Decoder3_212 (.dis(wire_438), .sel0(wire_136), .sel1(wire_21), .sel2(wire_329), .out0(wire_351), .out1(wire_173), .out2(wire_443), .out3(wire_233), .out4(wire_150), .out5(wire_417), .out6(wire_374), .out7(wire_391));
  TC_Splitter8 # (.UUID(64'd448586870420520821 ^ UUID)) Splitter8_213 (.in(wire_203), .out0(wire_136), .out1(wire_21), .out2(wire_329), .out3(wire_240), .out4(wire_95), .out5(wire_140), .out6(), .out7());
  TC_Or3 # (.UUID(64'd1235965720506732026 ^ UUID), .BIT_WIDTH(64'd1)) Or3_214 (.in0(wire_383), .in1(wire_41), .in2(wire_416), .out(wire_67));
  TC_Or3 # (.UUID(64'd64656781117703189 ^ UUID), .BIT_WIDTH(64'd1)) Or3_215 (.in0(wire_30[0:0]), .in1(wire_277), .in2(wire_86), .out(wire_458));
  TC_Not # (.UUID(64'd3756682246155706392 ^ UUID), .BIT_WIDTH(64'd1)) Not_216 (.in(wire_240), .out(wire_145));
  TC_Or3 # (.UUID(64'd1985979777212458751 ^ UUID), .BIT_WIDTH(64'd1)) Or3_217 (.in0(wire_61), .in1(wire_287[0:0]), .in2(wire_398), .out(wire_438));
  TC_Or3 # (.UUID(64'd1657864677517986892 ^ UUID), .BIT_WIDTH(64'd1)) Or3_218 (.in0(wire_51[0:0]), .in1(wire_113), .in2(wire_125), .out(wire_115));
  TC_And # (.UUID(64'd422870372255371239 ^ UUID), .BIT_WIDTH(64'd1)) And_219 (.in0(wire_145), .in1(wire_95), .out(wire_366));
  TC_Splitter8 # (.UUID(64'd760659632282220270 ^ UUID)) Splitter8_220 (.in(wire_130), .out0(wire_47), .out1(wire_155), .out2(wire_275), .out3(wire_277), .out4(wire_86), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd4082907615726159469 ^ UUID), .BIT_WIDTH(64'd1)) And_221 (.in0(wire_86), .in1(wire_216), .out(wire_461));
  TC_Splitter8 # (.UUID(64'd638362282452151696 ^ UUID)) Splitter8_222 (.in(wire_127), .out0(wire_244), .out1(wire_225), .out2(wire_74), .out3(wire_113), .out4(wire_125), .out5(), .out6(), .out7());
  TC_And # (.UUID(64'd3337535575473260291 ^ UUID), .BIT_WIDTH(64'd1)) And_223 (.in0(wire_125), .in1(wire_384), .out(wire_185));
  TC_Not # (.UUID(64'd558454314996824891 ^ UUID), .BIT_WIDTH(64'd1)) Not_224 (.in(wire_113), .out(wire_384));
  TC_Maker32 # (.UUID(64'd1972774908657050676 ^ UUID)) Maker32_225 (.in0(wire_202), .in1(wire_175), .in2(wire_129), .in3(wire_201), .out(wire_69));
  TC_Or # (.UUID(64'd2498810294022311638 ^ UUID), .BIT_WIDTH(64'd1)) Or_226 (.in0(wire_274), .in1(wire_296), .out(wire_105));
  TC_Switch # (.UUID(64'd2854933611415915645 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_227 (.en(wire_126), .in(wire_2), .out(wire_13_1[7:0]));
  TC_Or3 # (.UUID(64'd4211290242648182257 ^ UUID), .BIT_WIDTH(64'd1)) Or3_228 (.in0(wire_187), .in1(wire_89), .in2(wire_193), .out(wire_146));
  TC_Or # (.UUID(64'd4406510584467674262 ^ UUID), .BIT_WIDTH(64'd1)) Or_229 (.in0(wire_89), .in1(wire_193), .out(wire_61));
  TC_Or # (.UUID(64'd240802604651373700 ^ UUID), .BIT_WIDTH(64'd1)) Or_230 (.in0(wire_240), .in1(wire_95), .out(wire_398));
  TC_Switch # (.UUID(64'd2012067482831613303 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_231 (.en(wire_65), .in(wire_13[7:0]), .out(wire_55));
  TC_And # (.UUID(64'd647954593887269646 ^ UUID), .BIT_WIDTH(64'd1)) And_232 (.in0(wire_277), .in1(wire_86), .out(wire_200));
  TC_Splitter16 # (.UUID(64'd2940418270800807678 ^ UUID)) Splitter16_233 (.in(wire_156), .out0(wire_30), .out1(wire_51));
  TC_Maker16 # (.UUID(64'd4473516211661289785 ^ UUID)) Maker16_234 (.in0(wire_254), .in1({{7{1'b0}}, wire_4 }), .out(wire_156));
  TC_Or3 # (.UUID(64'd1738768736642702813 ^ UUID), .BIT_WIDTH(64'd1)) Or3_235 (.in0(wire_291), .in1(wire_102), .in2(wire_204), .out(wire_310));
  TC_Program # (.UUID(64'd145079491480902460 ^ UUID), .WORD_WIDTH(64'd8), .DEFAULT_FILE_NAME("Program_2036D0761E9DB3C.w8.bin"), .ARG_SIG("Program_2036D0761E9DB3C=%s")) Program_236 (.clk(clk), .rst(rst), .address({{8{1'b0}}, wire_139 }), .out0(wire_5), .out1(wire_106), .out2(wire_91), .out3(wire_414));
  TC_Maker8 # (.UUID(64'd1035456733302755062 ^ UUID)) Maker8_237 (.in0(wire_460), .in1(wire_259), .in2(wire_478), .in3(wire_426), .in4(wire_396), .in5(wire_157), .in6(wire_303), .in7(wire_471), .out(wire_298));
  TC_Maker8 # (.UUID(64'd2456434871637931222 ^ UUID)) Maker8_238 (.in0(wire_59), .in1(wire_437), .in2(wire_316), .in3(wire_463), .in4(wire_58), .in5(wire_264), .in6(wire_132), .in7(wire_255), .out(wire_350));
  TC_Maker8 # (.UUID(64'd3513223065136968424 ^ UUID)) Maker8_239 (.in0(wire_343), .in1(wire_385), .in2(wire_38), .in3(wire_16), .in4(wire_294), .in5(wire_352), .in6(wire_450), .in7(wire_278), .out(wire_42));
  TC_Maker8 # (.UUID(64'd1825601602491397740 ^ UUID)) Maker8_240 (.in0(wire_439), .in1(wire_400), .in2(wire_1), .in3(wire_441), .in4(wire_425), .in5(wire_362), .in6(wire_36), .in7(wire_137), .out(wire_77));
  TC_Maker8 # (.UUID(64'd1745865444850980894 ^ UUID)) Maker8_241 (.in0(wire_339), .in1(wire_325), .in2(wire_279), .in3(wire_368), .in4(wire_409), .in5(wire_457), .in6(wire_153), .in7(wire_470), .out(wire_149));
  TC_Decoder3 # (.UUID(64'd1376866551219367151 ^ UUID)) Decoder3_242 (.dis(wire_434), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_460), .out1(wire_259), .out2(wire_478), .out3(wire_426), .out4(wire_396), .out5(wire_157), .out6(wire_303), .out7(wire_471));
  TC_Not # (.UUID(64'd3892446360753336815 ^ UUID), .BIT_WIDTH(64'd1)) Not_243 (.in(wire_192), .out(wire_408));
  TC_And # (.UUID(64'd4179221552546912061 ^ UUID), .BIT_WIDTH(64'd1)) And_244 (.in0(wire_379), .in1(wire_191), .out(wire_11));
  TC_And3 # (.UUID(64'd2297715684806568026 ^ UUID), .BIT_WIDTH(64'd1)) And3_245 (.in0(wire_44), .in1(wire_468), .in2(wire_11), .out(wire_192));
  TC_And3 # (.UUID(64'd2633609611006090989 ^ UUID), .BIT_WIDTH(64'd1)) And3_246 (.in0(wire_70), .in1(wire_174), .in2(wire_107), .out(wire_141));
  TC_Not # (.UUID(64'd56970039485497802 ^ UUID), .BIT_WIDTH(64'd1)) Not_247 (.in(wire_174), .out(wire_468));
  TC_And3 # (.UUID(64'd157480515429222722 ^ UUID), .BIT_WIDTH(64'd1)) And3_248 (.in0(wire_44), .in1(wire_159), .in2(wire_333), .out(wire_183));
  TC_And # (.UUID(64'd1147743772323798401 ^ UUID), .BIT_WIDTH(64'd1)) And_249 (.in0(wire_24), .in1(wire_381), .out(wire_333));
  TC_And3 # (.UUID(64'd2961654373844858751 ^ UUID), .BIT_WIDTH(64'd1)) And3_250 (.in0(wire_378), .in1(wire_462), .in2(wire_101), .out(wire_120));
  TC_And # (.UUID(64'd1232556783305000021 ^ UUID), .BIT_WIDTH(64'd1)) And_251 (.in0(wire_24), .in1(wire_429), .out(wire_101));
  TC_And3 # (.UUID(64'd1620892037098951275 ^ UUID), .BIT_WIDTH(64'd1)) And3_252 (.in0(wire_44), .in1(wire_174), .in2(wire_9), .out(wire_369));
  TC_And # (.UUID(64'd1371408702773465615 ^ UUID), .BIT_WIDTH(64'd1)) And_253 (.in0(wire_435), .in1(wire_432), .out(wire_9));
  TC_And # (.UUID(64'd3049298419274804630 ^ UUID), .BIT_WIDTH(64'd1)) And_254 (.in0(wire_78), .in1(wire_32), .out(wire_107));
  TC_Not # (.UUID(64'd3896788527662292178 ^ UUID), .BIT_WIDTH(64'd1)) Not_255 (.in(wire_124), .out(wire_381));
  TC_Not # (.UUID(64'd2213138914507652729 ^ UUID), .BIT_WIDTH(64'd1)) Not_256 (.in(wire_174), .out(wire_159));
  TC_Not # (.UUID(64'd1715481119645584737 ^ UUID), .BIT_WIDTH(64'd1)) Not_257 (.in(wire_44), .out(wire_378));
  TC_Not # (.UUID(64'd2417925915142348864 ^ UUID), .BIT_WIDTH(64'd1)) Not_258 (.in(wire_124), .out(wire_429));
  TC_Not # (.UUID(64'd865647248024099255 ^ UUID), .BIT_WIDTH(64'd1)) Not_259 (.in(wire_174), .out(wire_462));
  TC_Not # (.UUID(64'd4459952580690051433 ^ UUID), .BIT_WIDTH(64'd1)) Not_260 (.in(wire_124), .out(wire_432));
  TC_Not # (.UUID(64'd3744757988884230908 ^ UUID), .BIT_WIDTH(64'd1)) Not_261 (.in(wire_24), .out(wire_435));
  TC_Not # (.UUID(64'd3181492288517670769 ^ UUID), .BIT_WIDTH(64'd1)) Not_262 (.in(wire_44), .out(wire_70));
  TC_Not # (.UUID(64'd4419382503653182595 ^ UUID), .BIT_WIDTH(64'd1)) Not_263 (.in(wire_124), .out(wire_32));
  TC_Not # (.UUID(64'd2505404667242823753 ^ UUID), .BIT_WIDTH(64'd1)) Not_264 (.in(wire_24), .out(wire_78));
  TC_Not # (.UUID(64'd650493536224126421 ^ UUID), .BIT_WIDTH(64'd1)) Not_265 (.in(wire_124), .out(wire_191));
  TC_Not # (.UUID(64'd1035715928482157684 ^ UUID), .BIT_WIDTH(64'd1)) Not_266 (.in(wire_24), .out(wire_379));
  TC_Not # (.UUID(64'd676402644750042592 ^ UUID), .BIT_WIDTH(64'd1)) Not_267 (.in(wire_183), .out(wire_434));
  TC_Not # (.UUID(64'd1922324152531657568 ^ UUID), .BIT_WIDTH(64'd1)) Not_268 (.in(wire_120), .out(wire_403));
  TC_Not # (.UUID(64'd3073651411181082508 ^ UUID), .BIT_WIDTH(64'd1)) Not_269 (.in(wire_369), .out(wire_365));
  TC_Not # (.UUID(64'd2629117106074357545 ^ UUID), .BIT_WIDTH(64'd1)) Not_270 (.in(wire_141), .out(wire_321));
  TC_Splitter8 # (.UUID(64'd1502652460628628447 ^ UUID)) Splitter8_271 (.in(wire_83), .out0(wire_99), .out1(wire_23), .out2(wire_45), .out3(wire_44), .out4(wire_174), .out5(wire_24), .out6(wire_124), .out7());
  TC_Decoder3 # (.UUID(64'd3968224955618952521 ^ UUID)) Decoder3_272 (.dis(wire_403), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_59), .out1(wire_437), .out2(wire_316), .out3(wire_463), .out4(wire_58), .out5(wire_264), .out6(wire_132), .out7(wire_255));
  TC_Decoder3 # (.UUID(64'd3094842192674468786 ^ UUID)) Decoder3_273 (.dis(wire_365), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_343), .out1(wire_385), .out2(wire_38), .out3(wire_16), .out4(wire_294), .out5(wire_352), .out6(wire_450), .out7(wire_278));
  TC_Decoder3 # (.UUID(64'd2218654558410367342 ^ UUID)) Decoder3_274 (.dis(wire_321), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_439), .out1(wire_400), .out2(wire_1), .out3(wire_441), .out4(wire_425), .out5(wire_362), .out6(wire_36), .out7(wire_137));
  TC_Decoder3 # (.UUID(64'd887192851734690171 ^ UUID)) Decoder3_275 (.dis(wire_408), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_339), .out1(wire_325), .out2(wire_279), .out3(wire_368), .out4(wire_409), .out5(wire_457), .out6(wire_153), .out7(wire_470));
  TC_Nor # (.UUID(64'd3866626421952475378 ^ UUID), .BIT_WIDTH(64'd1)) Nor_276 (.in0(wire_239), .in1(wire_140), .out(wire_222));
  TC_Maker8 # (.UUID(64'd4459904450968457517 ^ UUID)) Maker8_277 (.in0(wire_26), .in1(wire_236), .in2(wire_148), .in3(wire_382), .in4(wire_164), .in5(wire_227), .in6(wire_397), .in7(wire_332), .out(wire_418));
  TC_Not # (.UUID(64'd4215428181913493385 ^ UUID), .BIT_WIDTH(64'd1)) Not_278 (.in(wire_24), .out(wire_469));
  TC_Not # (.UUID(64'd4032471281002111157 ^ UUID), .BIT_WIDTH(64'd1)) Not_279 (.in(wire_124), .out(wire_177));
  TC_Decoder3 # (.UUID(64'd996120352387108425 ^ UUID)) Decoder3_280 (.dis(wire_330), .sel0(wire_99), .sel1(wire_23), .sel2(wire_45), .out0(wire_26), .out1(wire_236), .out2(wire_148), .out3(wire_382), .out4(wire_164), .out5(wire_227), .out6(wire_397), .out7(wire_332));
  TC_And3 # (.UUID(64'd1830606390080270525 ^ UUID), .BIT_WIDTH(64'd1)) And3_281 (.in0(wire_469), .in1(wire_177), .in2(wire_65), .out(wire_324));
  TC_Add # (.UUID(64'd4408145621911691017 ^ UUID), .BIT_WIDTH(64'd8)) Add8_282 (.in0(wire_288), .in1(wire_272), .ci(1'd0), .out(wire_83), .co());
  TC_Constant # (.UUID(64'd648021868671220940 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_283 (.out(wire_349));
  TC_Not # (.UUID(64'd4458448501919401293 ^ UUID), .BIT_WIDTH(64'd1)) Not_284 (.in(wire_44), .out(wire_241));
  TC_Not # (.UUID(64'd2656919742901693000 ^ UUID), .BIT_WIDTH(64'd1)) Not_285 (.in(wire_174), .out(wire_212));
  TC_Not # (.UUID(64'd1230714453098364340 ^ UUID), .BIT_WIDTH(64'd1)) Not_286 (.in(wire_289), .out(wire_330));
  TC_And3 # (.UUID(64'd1897262313226536408 ^ UUID), .BIT_WIDTH(64'd1)) And3_287 (.in0(wire_241), .in1(wire_212), .in2(wire_324), .out(wire_289));
  TC_Constant # (.UUID(64'd2443421582234399527 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h800000)) Constant32_288 (.out(wire_84));
  TC_And # (.UUID(64'd1571349306791071803 ^ UUID), .BIT_WIDTH(64'd8)) And8_289 (.in0(wire_363), .in1(wire_55), .out(wire_272));
  TC_Mux # (.UUID(64'd551248097054278276 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_290 (.sel(wire_134), .in0(wire_380), .in1(wire_360), .out(wire_76));
  TC_Constant # (.UUID(64'd3964982961058753694 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_291 (.out(wire_182));
  TC_Constant # (.UUID(64'd2589198461830330308 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h60)) Constant8_292 (.out(wire_388));
  TC_Constant # (.UUID(64'd2476831490286070788 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h30)) Constant8_293 (.out(wire_96));
  TC_Neg # (.UUID(64'd274447657020691882 ^ UUID), .BIT_WIDTH(64'd8)) Neg8_294 (.in(wire_284), .out(wire_288));
  TC_Switch # (.UUID(64'd4479910173006402860 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_295 (.en(wire_292), .in(wire_388), .out(wire_284_0));
  TC_Switch # (.UUID(64'd2036195697520703824 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_296 (.en(wire_355), .in(wire_96), .out(wire_284_1));
  TC_DotMatrixDisplay # (.UUID(64'd1118507987693416167 ^ UUID)) DotMatrixDisplay_297 (.clk(clk), .rst(rst), .en_y(wire_35[0:0]), .en_x(wire_76[0:0]), .color_info(wire_35), .pixel_info(wire_76));
  TC_DotMatrixDisplay # (.UUID(64'd1759213735214961697 ^ UUID)) DotMatrixDisplay_298 (.clk(clk), .rst(rst), .en_y(wire_31[0:0]), .en_x(wire_76[0:0]), .color_info(wire_31), .pixel_info(wire_76));
  TC_DotMatrixDisplay # (.UUID(64'd1992890972326438770 ^ UUID)) DotMatrixDisplay_299 (.clk(clk), .rst(rst), .en_y(wire_300[0:0]), .en_x(wire_76[0:0]), .color_info(wire_300), .pixel_info(wire_76));
  TC_Constant # (.UUID(64'd245597550392237676 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h30)) Constant8_300 (.out(wire_326));
  TC_Maker32 # (.UUID(64'd4070055319567765345 ^ UUID)) Maker32_301 (.in0({{7{1'b0}}, wire_163 }), .in1(wire_354), .in2(wire_476), .in3(wire_234), .out(wire_31));
  TC_LessU # (.UUID(64'd4201381607904528928 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_302 (.in0(wire_272), .in1(wire_421), .out(wire_165));
  TC_LessU # (.UUID(64'd1180503948796030951 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_303 (.in0(wire_272), .in1(wire_305), .out(wire_50));
  TC_LessU # (.UUID(64'd77917731117769392 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_304 (.in0(wire_272), .in1(wire_326), .out(wire_195));
  TC_Constant # (.UUID(64'd2240337880060160788 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h80)) Constant8_305 (.out(wire_421));
  TC_Constant # (.UUID(64'd4527172918742990571 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h60)) Constant8_306 (.out(wire_305));
  TC_Not # (.UUID(64'd778028366380114488 ^ UUID), .BIT_WIDTH(64'd1)) Not_307 (.in(wire_50), .out(wire_322));
  TC_Not # (.UUID(64'd4055431689765044358 ^ UUID), .BIT_WIDTH(64'd1)) Not_308 (.in(wire_195), .out(wire_8));
  TC_Not # (.UUID(64'd1010275238842509887 ^ UUID), .BIT_WIDTH(64'd1)) Not_309 (.in(wire_195), .out(wire_361));
  TC_And3 # (.UUID(64'd3539355440123382516 ^ UUID), .BIT_WIDTH(64'd1)) And3_310 (.in0(wire_8), .in1(wire_322), .in2(wire_165), .out(wire_292));
  TC_And3 # (.UUID(64'd3832948496576681869 ^ UUID), .BIT_WIDTH(64'd1)) And3_311 (.in0(wire_361), .in1(wire_50), .in2(wire_165), .out(wire_355));
  TC_And3 # (.UUID(64'd391397166249657057 ^ UUID), .BIT_WIDTH(64'd1)) And3_312 (.in0(wire_195), .in1(wire_50), .in2(wire_165), .out(wire_376));
  TC_Maker64 # (.UUID(64'd2613349598844013501 ^ UUID)) Maker64_313 (.in0({{7{1'b0}}, wire_349 }), .in1(wire_418), .in2(wire_149), .in3(wire_77), .in4(wire_42), .in5(wire_350), .in6(wire_298), .in7({{7{1'b0}}, wire_349 }), .out(wire_360));
  TC_Maker32 # (.UUID(64'd2223378423792437250 ^ UUID)) Maker32_314 (.in0({{7{1'b0}}, wire_81 }), .in1(wire_109), .in2(wire_268), .in3(wire_433), .out(wire_300));
  TC_Maker32 # (.UUID(64'd3989432137583600137 ^ UUID)) Maker32_315 (.in0({{7{1'b0}}, wire_110 }), .in1(wire_256), .in2(wire_473), .in3(wire_62), .out(wire_35));
  TC_Splitter32 # (.UUID(64'd505180353808894320 ^ UUID)) Splitter32_316 (.in(wire_114), .out0(), .out1(wire_256), .out2(wire_473), .out3(wire_62));
  TC_Splitter32 # (.UUID(64'd4136059224752756645 ^ UUID)) Splitter32_317 (.in(wire_114), .out0(), .out1(wire_354), .out2(wire_476), .out3(wire_234));
  TC_Splitter32 # (.UUID(64'd1271231891745783317 ^ UUID)) Splitter32_318 (.in(wire_114), .out0(), .out1(wire_109), .out2(wire_268), .out3(wire_433));
  TC_Constant # (.UUID(64'd3297416705186639367 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h1FFFFFFFFFFFF01)) Constant64_319 (.out(wire_308));
  TC_Mux # (.UUID(64'd1881013207545566499 ^ UUID), .BIT_WIDTH(64'd64)) Mux64_320 (.sel(wire_108), .in0(wire_308), .in1(wire_117), .out(wire_380));
  TC_Constant # (.UUID(64'd3348301751754001751 ^ UUID), .BIT_WIDTH(64'd64), .value(64'h10000FFFFFFFF01)) Constant64_321 (.out(wire_117));
  TC_Or # (.UUID(64'd2819938980275573952 ^ UUID), .BIT_WIDTH(64'd1)) Or_322 (.in0(wire_121), .in1(wire_292), .out(wire_81));
  TC_Or # (.UUID(64'd3147889042550481320 ^ UUID), .BIT_WIDTH(64'd1)) Or_323 (.in0(wire_309), .in1(wire_376), .out(wire_110));
  TC_DelayLine # (.UUID(64'd1341414154263104180 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_324 (.clk(clk), .rst(rst), .in(wire_197), .out(wire_271));
  TC_Constant # (.UUID(64'd1556929214979836766 ^ UUID), .BIT_WIDTH(64'd32), .value(32'h80000000)) Constant32_325 (.out(wire_64));
  TC_Switch # (.UUID(64'd3881038043152790915 ^ UUID), .BIT_WIDTH(64'd32)) Switch32_326 (.en(wire_222), .in(wire_84), .out(wire_248));
  TC_DelayLine # (.UUID(64'd2719614324323444454 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_327 (.clk(clk), .rst(rst), .in(wire_271), .out(wire_226));
  TC_Switch # (.UUID(64'd4603379206980955875 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_328 (.en(wire_239), .in(wire_271), .out(wire_121));
  TC_Not # (.UUID(64'd4292095226833103525 ^ UUID), .BIT_WIDTH(64'd1)) Not_329 (.in(wire_226), .out(wire_239));
  TC_Mux # (.UUID(64'd4236242586717471144 ^ UUID), .BIT_WIDTH(64'd32)) Mux32_330 (.sel(wire_286), .in0(wire_248), .in1(wire_64), .out(wire_114));
  TC_LessU # (.UUID(64'd3198049240392851104 ^ UUID), .BIT_WIDTH(64'd8)) LessU8_331 (.in0(wire_363), .in1(wire_55), .out(wire_286));
  TC_Constant # (.UUID(64'd1136323312820302173 ^ UUID), .BIT_WIDTH(64'd8), .value(8'h7F)) Constant8_332 (.out(wire_363));
  TC_Or # (.UUID(64'd3244493532244578566 ^ UUID), .BIT_WIDTH(64'd1)) Or_333 (.in0(wire_309), .in1(wire_355), .out(wire_163));
  TC_Switch # (.UUID(64'd1380797190081937409 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_334 (.en(wire_111), .in(wire_197), .out(wire_309));
  TC_Not # (.UUID(64'd4112928203054660527 ^ UUID), .BIT_WIDTH(64'd1)) Not_335 (.in(wire_269), .out(wire_111));
  TC_DelayLine # (.UUID(64'd3386030861920000876 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_336 (.clk(clk), .rst(rst), .in(wire_197), .out(wire_269));
  TC_Constant # (.UUID(64'd2747154628586710315 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_337 (.out(wire_197));
  TC_DelayLine # (.UUID(64'd4033780705460835019 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_338 (.clk(clk), .rst(rst), .in(wire_182), .out(wire_108));
  TC_DelayLine # (.UUID(64'd1957986231575802253 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_339 (.clk(clk), .rst(rst), .in(wire_108), .out(wire_134));
  TC_Timing # (.UUID(64'd191949461197767166 ^ UUID)) Timing_340 (.en(wire_472), .out(wire_122));
  TC_Not # (.UUID(64'd669353491571454392 ^ UUID), .BIT_WIDTH(64'd1)) Not_341 (.in(wire_131), .out(wire_243));
  TC_DelayLine # (.UUID(64'd3386813234232563563 ^ UUID), .BIT_WIDTH(64'd1)) DelayLine1_342 (.clk(clk), .rst(rst), .in(wire_427), .out(wire_131));
  TC_Switch # (.UUID(64'd1621668819963791229 ^ UUID), .BIT_WIDTH(64'd1)) Switch1_343 (.en(wire_243), .in(wire_54), .out(wire_427));
  TC_Or3 # (.UUID(64'd3441812953425143944 ^ UUID), .BIT_WIDTH(64'd1)) Or3_344 (.in0(wire_198[0:0]), .in1(wire_131), .in2(wire_209[0:0]), .out(wire_54));
  TC_Switch # (.UUID(64'd2666138502452780236 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_345 (.en(wire_198[0:0]), .in({{7{1'b0}}, wire_348 }), .out(wire_2_5));
  TC_Switch # (.UUID(64'd830658564569826705 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_346 (.en(wire_209[0:0]), .in({{7{1'b0}}, wire_348 }), .out(wire_0_5));
  TC_Constant # (.UUID(64'd3286728946413628039 ^ UUID), .BIT_WIDTH(64'd1), .value(1'd1)) On_347 (.out(wire_472));
  TC_Splitter16 # (.UUID(64'd1089016793051500988 ^ UUID)) Splitter16_348 (.in(wire_266), .out0(wire_209), .out1(wire_198));
  TC_Maker16 # (.UUID(64'd249508002051510401 ^ UUID)) Maker16_349 (.in0(wire_464), .in1(wire_430), .out(wire_266));
  TC_Splitter8 # (.UUID(64'd3424845306457333027 ^ UUID)) Splitter8_350 (.in(wire_299), .out0(), .out1(), .out2(wire_465), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Splitter64 # (.UUID(64'd196912585129497673 ^ UUID)) Splitter64_351 (.in(wire_122), .out0(), .out1(), .out2(wire_299), .out3(), .out4(), .out5(), .out6(), .out7());
  TC_Switch # (.UUID(64'd3742298234286761187 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_352 (.en(wire_304[0:0]), .in({{7{1'b0}}, wire_465 }), .out(wire_2_6));
  TC_Switch # (.UUID(64'd2409838377192211521 ^ UUID), .BIT_WIDTH(64'd8)) Switch8_353 (.en(wire_224[0:0]), .in(wire_122[7:0]), .out(wire_0_4));
  TC_Splitter32 # (.UUID(64'd118883049891919247 ^ UUID)) Splitter32_354 (.in(wire_359), .out0(wire_464), .out1(wire_430), .out2(wire_304), .out3(wire_224));
  TC_Maker32 # (.UUID(64'd301436605279209428 ^ UUID)) Maker32_355 (.in0({{7{1'b0}}, wire_200 }), .in1({{7{1'b0}}, wire_144 }), .in2({{7{1'b0}}, wire_27 }), .in3({{7{1'b0}}, wire_265 }), .out(wire_359));
  TC_Not # (.UUID(64'd2924370506823732469 ^ UUID), .BIT_WIDTH(64'd1)) Not_356 (.in(wire_277), .out(wire_480));
  TC_Not # (.UUID(64'd1358565458931546622 ^ UUID), .BIT_WIDTH(64'd1)) Not_357 (.in(wire_277), .out(wire_216));
  TC_Maker32 # (.UUID(64'd3731905900420244009 ^ UUID)) Maker32_358 (.in0({{7{1'b0}}, wire_112 }), .in1({{7{1'b0}}, wire_445 }), .in2({{7{1'b0}}, wire_452 }), .in3({{7{1'b0}}, wire_467 }), .out(wire_404));
  TC_Splitter32 # (.UUID(64'd3952628877771949754 ^ UUID)) Splitter32_359 (.in(wire_404), .out0(wire_158), .out1(wire_66), .out2(wire_261), .out3(wire_431));
  TC_Or # (.UUID(64'd1464181653386223728 ^ UUID), .BIT_WIDTH(64'd1)) Or_360 (.in0(wire_25), .in1(wire_68), .out(wire_186));
  TC_Or # (.UUID(64'd1071650078955089329 ^ UUID), .BIT_WIDTH(64'd1)) Or_361 (.in0(wire_345), .in1(wire_402), .out(wire_416));
  TC_Or # (.UUID(64'd3984947405899213483 ^ UUID), .BIT_WIDTH(64'd1)) Or_362 (.in0(wire_219), .in1(wire_229), .out(wire_143));
  TC_Or # (.UUID(64'd19590702580144813 ^ UUID), .BIT_WIDTH(64'd1)) Or_363 (.in0(wire_28), .in1(wire_211), .out(wire_442));
  TC_Decoder2 # (.UUID(64'd2363697850107914081 ^ UUID)) Decoder2_364 (.sel0(wire_431[0:0]), .sel1(wire_401), .out0(wire_449), .out1(wire_180), .out2(wire_474), .out3(wire_412));

  wire [7:0] wire_0;
  wire [7:0] wire_0_0;
  wire [7:0] wire_0_1;
  wire [7:0] wire_0_2;
  wire [7:0] wire_0_3;
  wire [7:0] wire_0_4;
  wire [7:0] wire_0_5;
  wire [7:0] wire_0_6;
  wire [7:0] wire_0_7;
  wire [7:0] wire_0_8;
  wire [7:0] wire_0_9;
  wire [7:0] wire_0_10;
  wire [7:0] wire_0_11;
  wire [7:0] wire_0_12;
  wire [7:0] wire_0_13;
  wire [7:0] wire_0_14;
  wire [7:0] wire_0_15;
  wire [7:0] wire_0_16;
  wire [7:0] wire_0_17;
  wire [7:0] wire_0_18;
  assign wire_0 = wire_0_0|wire_0_1|wire_0_2|wire_0_3|wire_0_4|wire_0_5|wire_0_6|wire_0_7|wire_0_8|wire_0_9|wire_0_10|wire_0_11|wire_0_12|wire_0_13|wire_0_14|wire_0_15|wire_0_16|wire_0_17|wire_0_18;
  wire [0:0] wire_1;
  wire [7:0] wire_2;
  wire [7:0] wire_2_0;
  wire [7:0] wire_2_1;
  wire [7:0] wire_2_2;
  wire [7:0] wire_2_3;
  wire [7:0] wire_2_4;
  wire [7:0] wire_2_5;
  wire [7:0] wire_2_6;
  wire [7:0] wire_2_7;
  wire [7:0] wire_2_8;
  wire [7:0] wire_2_9;
  wire [7:0] wire_2_10;
  wire [7:0] wire_2_11;
  wire [7:0] wire_2_12;
  wire [7:0] wire_2_13;
  wire [7:0] wire_2_14;
  wire [7:0] wire_2_15;
  wire [7:0] wire_2_16;
  wire [7:0] wire_2_17;
  wire [7:0] wire_2_18;
  assign wire_2 = wire_2_0|wire_2_1|wire_2_2|wire_2_3|wire_2_4|wire_2_5|wire_2_6|wire_2_7|wire_2_8|wire_2_9|wire_2_10|wire_2_11|wire_2_12|wire_2_13|wire_2_14|wire_2_15|wire_2_16|wire_2_17|wire_2_18;
  wire [0:0] wire_3;
  wire [0:0] wire_4;
  wire [63:0] wire_5;
  wire [0:0] wire_6;
  wire [0:0] wire_7;
  wire [0:0] wire_8;
  wire [0:0] wire_9;
  wire [7:0] wire_10;
  wire [0:0] wire_11;
  wire [7:0] wire_12;
  wire [63:0] wire_13;
  wire [63:0] wire_13_0;
  wire [63:0] wire_13_1;
  wire [63:0] wire_13_2;
  wire [63:0] wire_13_3;
  wire [63:0] wire_13_4;
  wire [63:0] wire_13_5;
  wire [63:0] wire_13_6;
  wire [63:0] wire_13_7;
  wire [63:0] wire_13_8;
  wire [63:0] wire_13_9;
  wire [63:0] wire_13_10;
  wire [63:0] wire_13_11;
  wire [63:0] wire_13_12;
  wire [63:0] wire_13_13;
  wire [63:0] wire_13_14;
  wire [63:0] wire_13_15;
  wire [63:0] wire_13_16;
  wire [63:0] wire_13_17;
  wire [63:0] wire_13_18;
  wire [63:0] wire_13_19;
  assign wire_13 = wire_13_0|wire_13_1|wire_13_2|wire_13_3|wire_13_4|wire_13_5|wire_13_6|wire_13_7|wire_13_8|wire_13_9|wire_13_10|wire_13_11|wire_13_12|wire_13_13|wire_13_14|wire_13_15|wire_13_16|wire_13_17|wire_13_18|wire_13_19;
  wire [0:0] wire_14;
  wire [7:0] wire_15;
  wire [0:0] wire_16;
  wire [7:0] wire_17;
  wire [0:0] wire_18;
  wire [7:0] wire_19;
  wire [0:0] wire_20;
  wire [0:0] wire_21;
  wire [0:0] wire_22;
  wire [0:0] wire_23;
  wire [0:0] wire_24;
  wire [0:0] wire_25;
  wire [0:0] wire_26;
  wire [0:0] wire_27;
  wire [0:0] wire_28;
  wire [0:0] wire_29;
  wire [7:0] wire_30;
  wire [31:0] wire_31;
  wire [0:0] wire_32;
  wire [0:0] wire_33;
  wire [7:0] wire_34;
  wire [7:0] wire_34_0;
  wire [7:0] wire_34_1;
  assign wire_34 = wire_34_0|wire_34_1;
  wire [31:0] wire_35;
  wire [0:0] wire_36;
  wire [7:0] wire_37;
  wire [0:0] wire_38;
  wire [0:0] wire_39;
  wire [0:0] wire_40;
  wire [0:0] wire_41;
  wire [7:0] wire_42;
  wire [7:0] wire_43;
  wire [0:0] wire_44;
  wire [0:0] wire_45;
  wire [7:0] wire_46;
  wire [0:0] wire_47;
  wire [0:0] wire_48;
  wire [0:0] wire_49;
  wire [0:0] wire_50;
  wire [7:0] wire_51;
  wire [0:0] wire_52;
  wire [0:0] wire_53;
  wire [0:0] wire_54;
  wire [7:0] wire_55;
  wire [0:0] wire_56;
  wire [7:0] wire_57;
  wire [0:0] wire_58;
  wire [0:0] wire_59;
  wire [0:0] wire_60;
  wire [0:0] wire_61;
  wire [7:0] wire_62;
  wire [7:0] wire_63;
  wire [31:0] wire_64;
  wire [0:0] wire_65;
  wire [7:0] wire_66;
  wire [0:0] wire_67;
  wire [0:0] wire_68;
  wire [31:0] wire_69;
  wire [0:0] wire_70;
  wire [0:0] wire_71;
  wire [0:0] wire_72;
  wire [0:0] wire_72_0;
  wire [0:0] wire_72_1;
  wire [0:0] wire_72_2;
  wire [0:0] wire_72_3;
  wire [0:0] wire_72_4;
  wire [0:0] wire_72_5;
  wire [0:0] wire_72_6;
  wire [0:0] wire_72_7;
  assign wire_72 = wire_72_0|wire_72_1|wire_72_2|wire_72_3|wire_72_4|wire_72_5|wire_72_6|wire_72_7;
  wire [0:0] wire_73;
  wire [0:0] wire_74;
  wire [0:0] wire_75;
  wire [63:0] wire_76;
  wire [7:0] wire_77;
  wire [0:0] wire_78;
  wire [0:0] wire_79;
  wire [7:0] wire_80;
  wire [7:0] wire_80_0;
  wire [7:0] wire_80_1;
  wire [7:0] wire_80_2;
  assign wire_80 = wire_80_0|wire_80_1|wire_80_2;
  wire [0:0] wire_81;
  wire [0:0] wire_82;
  wire [7:0] wire_83;
  wire [31:0] wire_84;
  wire [0:0] wire_85;
  wire [0:0] wire_86;
  wire [0:0] wire_87;
  wire [7:0] wire_88;
  wire [0:0] wire_89;
  wire [0:0] wire_90;
  wire [63:0] wire_91;
  wire [0:0] wire_92;
  wire [0:0] wire_93;
  wire [0:0] wire_94;
  wire [0:0] wire_95;
  wire [7:0] wire_96;
  wire [7:0] wire_97;
  wire [0:0] wire_98;
  wire [0:0] wire_99;
  wire [0:0] wire_100;
  wire [0:0] wire_101;
  wire [0:0] wire_102;
  wire [0:0] wire_103;
  wire [0:0] wire_104;
  wire [0:0] wire_105;
  wire [63:0] wire_106;
  wire [0:0] wire_107;
  wire [0:0] wire_108;
  wire [7:0] wire_109;
  wire [0:0] wire_110;
  wire [0:0] wire_111;
  wire [0:0] wire_112;
  wire [0:0] wire_113;
  wire [31:0] wire_114;
  wire [0:0] wire_115;
  wire [7:0] wire_116;
  wire [63:0] wire_117;
  wire [0:0] wire_118;
  wire [0:0] wire_119;
  wire [0:0] wire_120;
  wire [0:0] wire_121;
  wire [63:0] wire_122;
  wire [0:0] wire_123;
  wire [0:0] wire_124;
  wire [0:0] wire_125;
  wire [0:0] wire_126;
  wire [7:0] wire_127;
  wire [7:0] wire_128;
  wire [7:0] wire_128_0;
  wire [7:0] wire_128_1;
  assign wire_128 = wire_128_0|wire_128_1;
  wire [7:0] wire_129;
  wire [7:0] wire_130;
  wire [0:0] wire_131;
  wire [0:0] wire_132;
  wire [0:0] wire_133;
  wire [0:0] wire_134;
  wire [7:0] wire_135;
  wire [0:0] wire_136;
  wire [0:0] wire_137;
  wire [0:0] wire_138;
  wire [7:0] wire_139;
  wire [0:0] wire_140;
  wire [0:0] wire_141;
  wire [7:0] wire_142;
  wire [0:0] wire_143;
  wire [0:0] wire_144;
  wire [0:0] wire_145;
  wire [0:0] wire_146;
  wire [0:0] wire_147;
  wire [0:0] wire_148;
  wire [7:0] wire_149;
  wire [0:0] wire_150;
  wire [0:0] wire_151;
  wire [7:0] wire_152;
  wire [0:0] wire_153;
  wire [0:0] wire_154;
  wire [0:0] wire_155;
  wire [15:0] wire_156;
  wire [0:0] wire_157;
  wire [7:0] wire_158;
  wire [0:0] wire_159;
  wire [7:0] wire_160;
  wire [7:0] wire_161;
  wire [0:0] wire_162;
  wire [0:0] wire_163;
  wire [0:0] wire_164;
  wire [0:0] wire_165;
  wire [0:0] wire_166;
  wire [7:0] wire_167;
  wire [7:0] wire_168;
  wire [7:0] wire_168_0;
  wire [7:0] wire_168_1;
  assign wire_168 = wire_168_0|wire_168_1;
  wire [0:0] wire_169;
  wire [0:0] wire_170;
  wire [0:0] wire_171;
  wire [0:0] wire_172;
  wire [0:0] wire_173;
  wire [0:0] wire_174;
  wire [7:0] wire_175;
  wire [0:0] wire_176;
  wire [0:0] wire_177;
  wire [0:0] wire_178;
  wire [0:0] wire_179;
  wire [0:0] wire_180;
  wire [63:0] wire_181;
  wire [0:0] wire_182;
  wire [0:0] wire_183;
  wire [0:0] wire_184;
  wire [0:0] wire_185;
  wire [0:0] wire_186;
  wire [0:0] wire_187;
  wire [0:0] wire_188;
  wire [7:0] wire_189;
  wire [7:0] wire_190;
  wire [0:0] wire_191;
  wire [0:0] wire_192;
  wire [0:0] wire_193;
  wire [0:0] wire_194;
  wire [0:0] wire_195;
  wire [0:0] wire_196;
  wire [0:0] wire_197;
  wire [7:0] wire_198;
  wire [0:0] wire_199;
  wire [0:0] wire_200;
  wire [7:0] wire_201;
  wire [7:0] wire_202;
  wire [7:0] wire_203;
  wire [0:0] wire_204;
  wire [0:0] wire_205;
  wire [0:0] wire_206;
  wire [0:0] wire_207;
  wire [7:0] wire_208;
  wire [7:0] wire_209;
  wire [0:0] wire_210;
  wire [0:0] wire_211;
  wire [0:0] wire_212;
  wire [0:0] wire_213;
  wire [15:0] wire_214;
  wire [7:0] wire_215;
  wire [7:0] wire_215_0;
  wire [7:0] wire_215_1;
  assign wire_215 = wire_215_0|wire_215_1;
  wire [0:0] wire_216;
  wire [0:0] wire_217;
  wire [0:0] wire_218;
  wire [0:0] wire_219;
  wire [0:0] wire_220;
  wire [0:0] wire_221;
  wire [0:0] wire_222;
  wire [0:0] wire_223;
  wire [7:0] wire_224;
  wire [0:0] wire_225;
  wire [0:0] wire_226;
  wire [0:0] wire_227;
  wire [0:0] wire_228;
  wire [0:0] wire_229;
  wire [7:0] wire_230;
  wire [7:0] wire_231;
  wire [0:0] wire_232;
  wire [0:0] wire_233;
  wire [7:0] wire_234;
  wire [0:0] wire_235;
  wire [0:0] wire_236;
  wire [7:0] wire_237;
  wire [7:0] wire_238;
  wire [0:0] wire_239;
  wire [0:0] wire_240;
  wire [0:0] wire_241;
  wire [0:0] wire_242;
  wire [0:0] wire_243;
  wire [0:0] wire_244;
  wire [0:0] wire_245;
  wire [0:0] wire_246;
  wire [0:0] wire_247;
  wire [31:0] wire_248;
  wire [0:0] wire_249;
  wire [0:0] wire_250;
  wire [0:0] wire_251;
  wire [7:0] wire_252;
  wire [0:0] wire_253;
  wire [7:0] wire_254;
  wire [0:0] wire_255;
  wire [7:0] wire_256;
  wire [0:0] wire_257;
  wire [7:0] wire_258;
  wire [0:0] wire_259;
  wire [7:0] wire_260;
  wire [7:0] wire_261;
  wire [0:0] wire_262;
  wire [0:0] wire_263;
  wire [0:0] wire_264;
  wire [0:0] wire_265;
  wire [15:0] wire_266;
  wire [0:0] wire_267;
  wire [7:0] wire_268;
  wire [0:0] wire_269;
  wire [7:0] wire_270;
  wire [0:0] wire_271;
  wire [7:0] wire_272;
  wire [7:0] wire_273;
  wire [0:0] wire_274;
  wire [0:0] wire_275;
  wire [0:0] wire_276;
  wire [0:0] wire_277;
  wire [0:0] wire_278;
  wire [0:0] wire_279;
  wire [7:0] wire_280;
  wire [0:0] wire_281;
  wire [7:0] wire_282;
  wire [7:0] wire_283;
  wire [7:0] wire_284;
  wire [7:0] wire_284_0;
  wire [7:0] wire_284_1;
  assign wire_284 = wire_284_0|wire_284_1;
  wire [0:0] wire_285;
  wire [0:0] wire_286;
  wire [7:0] wire_287;
  wire [7:0] wire_288;
  wire [0:0] wire_289;
  wire [0:0] wire_290;
  wire [0:0] wire_291;
  wire [0:0] wire_292;
  wire [0:0] wire_293;
  wire [0:0] wire_294;
  wire [7:0] wire_295;
  wire [0:0] wire_296;
  wire [7:0] wire_297;
  wire [7:0] wire_297_0;
  wire [7:0] wire_297_1;
  assign wire_297 = wire_297_0|wire_297_1;
  wire [7:0] wire_298;
  wire [7:0] wire_299;
  wire [31:0] wire_300;
  wire [0:0] wire_301;
  wire [0:0] wire_302;
  wire [0:0] wire_303;
  wire [7:0] wire_304;
  wire [7:0] wire_305;
  wire [0:0] wire_306;
  wire [0:0] wire_307;
  wire [63:0] wire_308;
  wire [0:0] wire_309;
  wire [0:0] wire_310;
  wire [7:0] wire_311;
  wire [7:0] wire_312;
  wire [7:0] wire_313;
  wire [0:0] wire_314;
  wire [0:0] wire_315;
  wire [0:0] wire_316;
  wire [7:0] wire_317;
  wire [0:0] wire_318;
  wire [7:0] wire_319;
  wire [0:0] wire_320;
  wire [0:0] wire_321;
  wire [0:0] wire_322;
  wire [7:0] wire_323;
  wire [0:0] wire_324;
  wire [0:0] wire_325;
  wire [7:0] wire_326;
  wire [7:0] wire_327;
  wire [7:0] wire_328;
  wire [0:0] wire_329;
  wire [0:0] wire_330;
  wire [0:0] wire_331;
  wire [0:0] wire_332;
  wire [0:0] wire_333;
  wire [0:0] wire_334;
  wire [0:0] wire_335;
  wire [0:0] wire_336;
  wire [0:0] wire_337;
  wire [0:0] wire_338;
  wire [0:0] wire_339;
  wire [7:0] wire_340;
  wire [0:0] wire_341;
  wire [0:0] wire_342;
  wire [0:0] wire_343;
  wire [15:0] wire_344;
  wire [0:0] wire_345;
  wire [7:0] wire_346;
  wire [0:0] wire_347;
  wire [0:0] wire_348;
  assign wire_348 = 0;
  wire [0:0] wire_349;
  wire [7:0] wire_350;
  wire [0:0] wire_351;
  wire [0:0] wire_352;
  wire [0:0] wire_353;
  wire [7:0] wire_354;
  wire [0:0] wire_355;
  wire [7:0] wire_356;
  wire [15:0] wire_357;
  wire [7:0] wire_358;
  wire [31:0] wire_359;
  wire [63:0] wire_360;
  wire [0:0] wire_361;
  wire [0:0] wire_362;
  wire [7:0] wire_363;
  wire [7:0] wire_364;
  wire [0:0] wire_365;
  wire [0:0] wire_366;
  wire [7:0] wire_367;
  wire [0:0] wire_368;
  wire [0:0] wire_369;
  wire [0:0] wire_370;
  wire [0:0] wire_371;
  wire [0:0] wire_372;
  wire [0:0] wire_373;
  wire [0:0] wire_374;
  wire [0:0] wire_375;
  wire [0:0] wire_376;
  wire [0:0] wire_377;
  wire [0:0] wire_378;
  wire [0:0] wire_379;
  wire [63:0] wire_380;
  wire [0:0] wire_381;
  wire [0:0] wire_382;
  wire [0:0] wire_383;
  wire [0:0] wire_384;
  wire [0:0] wire_385;
  wire [7:0] wire_386;
  wire [0:0] wire_387;
  wire [7:0] wire_388;
  wire [7:0] wire_389;
  wire [0:0] wire_390;
  wire [0:0] wire_391;
  wire [7:0] wire_392;
  wire [0:0] wire_393;
  assign wire_393 = 0;
  wire [0:0] wire_394;
  wire [0:0] wire_395;
  wire [0:0] wire_396;
  wire [0:0] wire_397;
  wire [0:0] wire_398;
  wire [7:0] wire_399;
  wire [0:0] wire_400;
  wire [0:0] wire_401;
  wire [0:0] wire_402;
  wire [0:0] wire_403;
  wire [31:0] wire_404;
  wire [0:0] wire_405;
  wire [7:0] wire_406;
  wire [0:0] wire_407;
  wire [0:0] wire_408;
  wire [0:0] wire_409;
  wire [0:0] wire_410;
  wire [7:0] wire_411;
  wire [0:0] wire_412;
  wire [0:0] wire_413;
  wire [63:0] wire_414;
  wire [7:0] wire_415;
  wire [0:0] wire_416;
  wire [0:0] wire_417;
  wire [7:0] wire_418;
  wire [0:0] wire_419;
  wire [0:0] wire_420;
  wire [7:0] wire_421;
  wire [0:0] wire_422;
  wire [0:0] wire_423;
  wire [7:0] wire_424;
  wire [0:0] wire_425;
  wire [0:0] wire_426;
  wire [0:0] wire_427;
  wire [7:0] wire_428;
  wire [0:0] wire_429;
  wire [7:0] wire_430;
  wire [7:0] wire_431;
  wire [0:0] wire_432;
  wire [7:0] wire_433;
  wire [0:0] wire_434;
  wire [0:0] wire_435;
  wire [7:0] wire_436;
  wire [0:0] wire_437;
  wire [0:0] wire_438;
  wire [0:0] wire_439;
  wire [0:0] wire_440;
  wire [0:0] wire_441;
  wire [0:0] wire_442;
  wire [0:0] wire_443;
  wire [0:0] wire_444;
  wire [0:0] wire_445;
  wire [7:0] wire_446;
  wire [0:0] wire_447;
  wire [7:0] wire_448;
  wire [0:0] wire_449;
  wire [0:0] wire_450;
  wire [0:0] wire_451;
  wire [0:0] wire_452;
  wire [7:0] wire_453;
  wire [0:0] wire_454;
  wire [0:0] wire_455;
  wire [7:0] wire_456;
  wire [0:0] wire_457;
  wire [0:0] wire_458;
  wire [0:0] wire_459;
  wire [0:0] wire_460;
  wire [0:0] wire_461;
  wire [0:0] wire_462;
  wire [0:0] wire_463;
  wire [7:0] wire_464;
  wire [0:0] wire_465;
  wire [7:0] wire_466;
  wire [0:0] wire_467;
  wire [0:0] wire_468;
  wire [0:0] wire_469;
  wire [0:0] wire_470;
  wire [0:0] wire_471;
  wire [0:0] wire_472;
  wire [7:0] wire_473;
  wire [0:0] wire_474;
  wire [7:0] wire_475;
  wire [7:0] wire_476;
  wire [7:0] wire_477;
  wire [0:0] wire_478;
  wire [7:0] wire_479;
  wire [0:0] wire_480;

endmodule
